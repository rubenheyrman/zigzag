//Hier for 'I_wr_data_rsci_idat_bfwt'
module temp_odc_impl_1451 ( I_wr_data_rsci_ivld_bfwt_0 , reg_I_wr_data_rsci_irdy_run_psct_cse_1
 , run_wten_2 , I_wr_data_rsci_bcwt_3 , I_mac_pntr_sva_4 , I_data_vld_sva_dfm_1_1_5
 , reg_W_instr_in_rsci_oswt_cse_1_6 , O_instr_in_rsci_bcwt_7 , I_instr_in_rsci_bcwt_8
 , W_instr_in_rsci_bcwt_9 , main_stage_0_2_10 , I_wr_pntr_sva_11 , state_var_12
 , O_instr_L1_out_rsci_bcwt_13 , reg_I_instr_L1_out_rsci_ivld_run_psct_cse_14
 , I_instr_L1_out_rsci_bcwt_15 , reg_W_instr_L1_out_rsci_ivld_run_psct_cse_16
 , W_instr_L1_out_rsci_bcwt_17 , reg_O_instr_L1_out_rsci_ivld_run_psct_cse_18
 , t_out ) ;
 input wire  I_wr_data_rsci_ivld_bfwt_0 ; 
 input wire  reg_I_wr_data_rsci_irdy_run_psct_cse_1 ; 
 input wire  run_wten_2 ; 
 input wire  I_wr_data_rsci_bcwt_3 ; 
 input wire  [4:0]  I_mac_pntr_sva_4 ; 
 input wire  I_data_vld_sva_dfm_1_1_5 ; 
 input wire  reg_W_instr_in_rsci_oswt_cse_1_6 ; 
 input wire  O_instr_in_rsci_bcwt_7 ; 
 input wire  I_instr_in_rsci_bcwt_8 ; 
 input wire  W_instr_in_rsci_bcwt_9 ; 
 input wire  main_stage_0_2_10 ; 
 input wire  [4:0]  I_wr_pntr_sva_11 ; 
 input wire  [0:0]  state_var_12 ; 
 input wire  O_instr_L1_out_rsci_bcwt_13 ; 
 input wire  reg_I_instr_L1_out_rsci_ivld_run_psct_cse_14 ; 
 input wire  I_instr_L1_out_rsci_bcwt_15 ; 
 input wire  reg_W_instr_L1_out_rsci_ivld_run_psct_cse_16 ; 
 input wire  W_instr_L1_out_rsci_bcwt_17 ; 
 input wire  reg_O_instr_L1_out_rsci_ivld_run_psct_cse_18 ; 
 output wire  t_out ; 
 wire E_273901 ; 
assign t_out = E_273901 ;
 wire E_273900 ; 
 wire E_273899 ; 
 wire E_273898 ; 
 wire E_273897 ; 
 wire E_273896 ; 
 wire E_273895 ; 
 wire E_273894 ; 
 wire E_273893 ; 
 wire E_273892 ; 
 wire E_273891 ; 
 wire E_273890 ; 
 wire E_273889 ; 
 wire E_273888 ; 
 wire E_273887 ; 
 wire E_273886 ; 
 wire E_273885 ; 
 wire E_273884 ; 
 wire E_273883 ; 
 wire E_273882 ; 
 wire E_273881 ; 
 wire E_273880 ; 
 wire E_273879 ; 
 wire E_273878 ; 
 wire E_273877 ; 
 wire E_273876 ; 
 wire E_273875 ; 
 wire E_273874 ; 
 wire E_273873 ; 
 wire E_273872 ; 
 wire E_273871 ; 
 wire E_273870 ; 
 wire E_273869 ; 
 wire E_273868 ; 
 wire E_273867 ; 
 wire E_273866 ; 
 wire E_273865 ; 
 wire E_273864 ; 
 wire E_273863 ; 
 wire E_273862 ; 
 wire E_273861 ; 
 wire E_273860 ; 
 wire E_273859 ; 
 wire E_273858 ; 
 wire E_273857 ; 
 wire E_273856 ; 
 wire E_273855 ; 
 wire E_273854 ; 
 wire E_273853 ; 
 wire E_273852 ; 
 wire E_273851 ; 
 wire E_273850 ; 
 wire E_273849 ; 
 wire E_273848 ; 
 wire E_273847 ; 
 wire E_273846 ; 
 wire E_273845 ; 
 wire E_273844 ; 
 wire E_273843 ; 
 wire E_273842 ; 
 wire E_273841 ; 
 wire E_273840 ; 
 wire E_273839 ; 
 wire E_273838 ; 
 wire E_273837 ; 
 wire E_273836 ; 
 wire E_273835 ; 
 wire E_273834 ; 
 wire E_273833 ; 
 wire E_273832 ; 
 wire E_273831 ; 
 wire E_273830 ; 
 wire E_273829 ; 
 wire E_273828 ; 
 wire E_273827 ; 
 wire E_273826 ; 
 wire E_273825 ; 
 wire E_273824 ; 
 wire E_273823 ; 
 wire E_273822 ; 
 wire E_273821 ; 
 wire E_273820 ; 
 wire E_273819 ; 
 wire E_273818 ; 
 wire E_273817 ; 
 wire E_273816 ; 
 wire E_273815 ; 
 wire E_273814 ; 
 wire E_273813 ; 
 wire E_273812 ; 
 wire E_273811 ; 
 wire E_273810 ; 
 wire E_273809 ; 
 wire E_273808 ; 
 wire E_273807 ; 
 wire E_273806 ; 
 wire E_273805 ; 
 wire E_273804 ; 
 wire E_273803 ; 
 wire E_273802 ; 
 wire E_273801 ; 
 wire E_273800 ; 
 wire E_273799 ; 
 wire E_273798 ; 
 wire E_273797 ; 
 wire E_273796 ; 
 wire E_273795 ; 
 wire E_273794 ; 
 wire E_273793 ; 
 wire E_273792 ; 
 wire E_273791 ; 
 wire E_273790 ; 
 wire E_273789 ; 
 wire E_273788 ; 
 wire E_273787 ; 
 wire E_273786 ; 
 wire E_273785 ; 
 wire E_273784 ; 
assign E_273784 = reg_O_instr_L1_out_rsci_ivld_run_psct_cse_18 ;
 wire E_273783 ; 
 wire E_273782 ; 
 wire E_273781 ; 
 wire E_273780 ; 
 wire E_273779 ; 
 wire E_273778 ; 
 wire E_273777 ; 
 wire E_273776 ; 
 wire E_273775 ; 
 wire E_273774 ; 
 wire E_273773 ; 
 wire E_273772 ; 
 wire E_273771 ; 
 wire E_273770 ; 
 wire E_273769 ; 
 wire E_273768 ; 
 wire E_273767 ; 
 wire E_273766 ; 
 wire E_273765 ; 
 wire E_273764 ; 
 wire E_273763 ; 
 wire E_273762 ; 
 wire E_273761 ; 
 wire E_273760 ; 
 wire E_273759 ; 
 wire E_273758 ; 
 wire E_273757 ; 
 wire E_273756 ; 
 wire E_273755 ; 
 wire E_273754 ; 
 wire E_273753 ; 
 wire E_273752 ; 
 wire E_273751 ; 
 wire E_273750 ; 
 wire E_273749 ; 
 wire E_273748 ; 
 wire E_273747 ; 
 wire E_273746 ; 
 wire E_273745 ; 
 wire E_273744 ; 
 wire E_273743 ; 
 wire E_273742 ; 
 wire E_273741 ; 
 wire E_273740 ; 
 wire E_273739 ; 
 wire E_273738 ; 
 wire E_273737 ; 
 wire E_273736 ; 
assign E_273736 = W_instr_L1_out_rsci_bcwt_17 ;
 wire E_273735 ; 
 wire E_273734 ; 
 wire E_273733 ; 
assign E_273733 = reg_W_instr_L1_out_rsci_ivld_run_psct_cse_16 ;
 wire E_273732 ; 
 wire E_273731 ; 
 wire E_273730 ; 
assign E_273730 = I_instr_L1_out_rsci_bcwt_15 ;
 wire E_273729 ; 
 wire E_273728 ; 
 wire E_273727 ; 
assign E_273727 = reg_I_instr_L1_out_rsci_ivld_run_psct_cse_14 ;
 wire E_273726 ; 
 wire E_273725 ; 
 wire E_273724 ; 
 wire E_273723 ; 
assign E_273723 = O_instr_L1_out_rsci_bcwt_13 ;
 wire E_273722 ; 
 wire E_273721 ; 
 wire E_273720 ; 
 wire E_273719 ; 
 wire E_273718 ; 
 wire E_273717 ; 
 wire E_273716 ; 
 wire E_273715 ; 
 wire E_273714 ; 
 wire E_273713 ; 
 wire E_273712 ; 
 wire E_273711 ; 
 wire E_273710 ; 
 wire E_273709 ; 
 wire E_273708 ; 
 wire E_273707 ; 
 wire E_273706 ; 
 wire E_273705 ; 
 wire E_273704 ; 
 wire E_273703 ; 
 wire E_273702 ; 
 wire E_273701 ; 
 wire E_273700 ; 
 wire E_273699 ; 
 wire E_273698 ; 
 wire E_273697 ; 
 wire E_273696 ; 
 wire E_273695 ; 
 wire E_273694 ; 
 wire E_273693 ; 
 wire E_273692 ; 
 wire E_273691 ; 
 wire E_273690 ; 
 wire E_273689 ; 
 wire E_273688 ; 
 wire E_273687 ; 
 wire E_273686 ; 
 wire E_273685 ; 
 wire E_273684 ; 
 wire E_273683 ; 
 wire E_273682 ; 
 wire E_273681 ; 
 wire E_273680 ; 
 wire E_273679 ; 
 wire E_273678 ; 
 wire E_273677 ; 
 wire E_273676 ; 
 wire E_273675 ; 
 wire E_273674 ; 
 wire E_273673 ; 
 wire E_273672 ; 
 wire E_273671 ; 
 wire E_273670 ; 
 wire E_273669 ; 
 wire E_273668 ; 
 wire E_273667 ; 
 wire E_273666 ; 
 wire E_273665 ; 
 wire E_273664 ; 
 wire E_273663 ; 
 wire E_273662 ; 
 wire E_273661 ; 
 wire E_273660 ; 
 wire E_273659 ; 
 wire E_273658 ; 
 wire E_273657 ; 
 wire E_273656 ; 
 wire E_273655 ; 
 wire E_273654 ; 
 wire E_273653 ; 
 wire E_273652 ; 
 wire E_273651 ; 
 wire E_273650 ; 
 wire E_273649 ; 
 wire E_273648 ; 
 wire E_273647 ; 
 wire E_273646 ; 
 wire E_273645 ; 
 wire E_273644 ; 
 wire E_273643 ; 
 wire  [0:0] E_273642 ; 
assign E_273642 = state_var_12 ;
 wire E_273641 ; 
 wire E_273640 ; 
 wire E_273639 ; 
 wire E_273638 ; 
 wire E_273637 ; 
 wire E_273636 ; 
 wire E_273635 ; 
 wire E_273634 ; 
 wire E_273633 ; 
 wire E_273632 ; 
 wire E_273631 ; 
 wire E_273630 ; 
 wire E_273629 ; 
 wire  [4:0] E_273628 ; 
assign E_273628 = I_wr_pntr_sva_11 ;
 wire E_273627 ; 
 wire E_273626 ; 
 wire E_273625 ; 
 wire E_273624 ; 
assign E_273624 = main_stage_0_2_10 ;
 wire E_273623 ; 
 wire E_273622 ; 
 wire E_273621 ; 
assign E_273621 = W_instr_in_rsci_bcwt_9 ;
 wire E_273620 ; 
 wire E_273619 ; 
assign E_273619 = I_instr_in_rsci_bcwt_8 ;
 wire E_273618 ; 
 wire E_273617 ; 
assign E_273617 = O_instr_in_rsci_bcwt_7 ;
 wire E_273616 ; 
 wire E_273615 ; 
 wire E_273614 ; 
assign E_273614 = reg_W_instr_in_rsci_oswt_cse_1_6 ;
 wire E_273613 ; 
 wire E_273612 ; 
 wire E_273611 ; 
 wire E_273610 ; 
 wire E_273609 ; 
 wire E_273608 ; 
 wire E_273607 ; 
 wire E_273606 ; 
 wire E_273605 ; 
 wire E_273604 ; 
assign E_273604 = I_data_vld_sva_dfm_1_1_5 ;
 wire E_273603 ; 
 wire E_273602 ; 
 wire E_273601 ; 
 wire E_273600 ; 
 wire E_273599 ; 
 wire E_273598 ; 
 wire E_273597 ; 
 wire E_273596 ; 
 wire E_273595 ; 
 wire E_273594 ; 
 wire E_273593 ; 
 wire E_273592 ; 
 wire E_273591 ; 
 wire E_273590 ; 
 wire  [4:0] E_273589 ; 
assign E_273589 = I_mac_pntr_sva_4 ;
 wire E_273588 ; 
 wire E_273587 ; 
 wire E_273586 ; 
 wire E_273585 ; 
 wire E_273584 ; 
assign E_273584 = I_wr_data_rsci_bcwt_3 ;
 wire E_273583 ; 
 wire E_273582 ; 
 wire E_273581 ; 
 wire E_273580 ; 
 wire E_273579 ; 
 wire E_273578 ; 
 wire E_273577 ; 
 wire E_273576 ; 
 wire E_273575 ; 
 wire E_273574 ; 
 wire E_273573 ; 
 wire E_273572 ; 
 wire E_273571 ; 
 wire E_273570 ; 
 wire E_273569 ; 
 wire E_273568 ; 
 wire E_273567 ; 
 wire E_273566 ; 
 wire E_273565 ; 
 wire E_273564 ; 
 wire E_273563 ; 
 wire E_273562 ; 
 wire E_273561 ; 
 wire E_273560 ; 
 wire E_273559 ; 
 wire E_273558 ; 
 wire E_273557 ; 
 wire E_273556 ; 
 wire E_273555 ; 
 wire E_273554 ; 
 wire E_273553 ; 
 wire E_273552 ; 
 wire E_273551 ; 
 wire E_273550 ; 
 wire E_273549 ; 
 wire E_273548 ; 
 wire E_273547 ; 
 wire E_273546 ; 
 wire E_273545 ; 
 wire E_273544 ; 
 wire E_273543 ; 
 wire E_273542 ; 
 wire E_273541 ; 
 wire E_273540 ; 
 wire E_273539 ; 
 wire E_273538 ; 
 wire E_273537 ; 
 wire E_273536 ; 
 wire E_273535 ; 
 wire E_273534 ; 
 wire E_273533 ; 
 wire E_273532 ; 
 wire E_273531 ; 
 wire E_273530 ; 
 wire E_273529 ; 
 wire E_273528 ; 
 wire E_273527 ; 
 wire E_273526 ; 
 wire E_273525 ; 
 wire E_273524 ; 
 wire E_273523 ; 
 wire E_273522 ; 
 wire E_273521 ; 
 wire E_273520 ; 
 wire E_273519 ; 
 wire E_273518 ; 
 wire E_273517 ; 
 wire E_273516 ; 
 wire E_273515 ; 
 wire E_273514 ; 
 wire E_273513 ; 
 wire E_273512 ; 
 wire E_273511 ; 
 wire E_273510 ; 
 wire E_273509 ; 
 wire E_273508 ; 
 wire E_273507 ; 
 wire E_273506 ; 
 wire E_273505 ; 
 wire E_273504 ; 
 wire E_273503 ; 
assign E_273503 = run_wten_2 ;
 wire E_273502 ; 
 wire E_273501 ; 
 wire E_273500 ; 
assign E_273500 = reg_I_wr_data_rsci_irdy_run_psct_cse_1 ;
 wire E_273499 ; 
 wire E_273498 ; 
assign E_273498 = I_wr_data_rsci_ivld_bfwt_0 ;
 wire E_273497 ; 
 wire E_273496 ; 
  assign /* unsigned    bit */  E_273901 = ( !E_273496 ) ;
  assign /* unsigned    bit */  E_273900 = (E_273588 & E_273740) ;
  assign /* unsigned    bit */  E_273899 = (E_273592 & E_273741) ;
  assign /* unsigned    bit */  E_273898 = (E_273595 & E_273742) ;
  assign /* unsigned    bit */  E_273897 = (E_273598 & E_273743) ;
  assign /* unsigned    bit */  E_273896 = (E_273601 & E_273744) ;
  assign /* unsigned    bit */  E_273895 = (E_273604 & E_273745) ;
  assign /* unsigned    bit */  E_273894 = (E_273588 & E_273797) ;
  assign /* unsigned    bit */  E_273893 = (E_273592 & E_273798) ;
  assign /* unsigned    bit */  E_273892 = (E_273595 & E_273799) ;
  assign /* unsigned    bit */  E_273891 = (E_273598 & E_273800) ;
  assign /* unsigned    bit */  E_273890 = (E_273601 & E_273801) ;
  assign /* unsigned    bit */  E_273889 = (E_273604 & E_273802) ;
  assign /* unsigned    bit */  E_273888 = (E_273588 & E_273774) ;
  assign /* unsigned    bit */  E_273887 = (E_273592 & E_273775) ;
  assign /* unsigned    bit */  E_273886 = (E_273595 & E_273776) ;
  assign /* unsigned    bit */  E_273885 = (E_273598 & E_273777) ;
  assign /* unsigned    bit */  E_273884 = (E_273601 & E_273778) ;
  assign /* unsigned    bit */  E_273883 = (E_273604 & E_273779) ;
  assign /* unsigned    bit */  E_273882 = (E_273588 & E_273829) ;
  assign /* unsigned    bit */  E_273881 = (E_273592 & E_273830) ;
  assign /* unsigned    bit */  E_273880 = (E_273595 & E_273831) ;
  assign /* unsigned    bit */  E_273879 = (E_273598 & E_273832) ;
  assign /* unsigned    bit */  E_273878 = (E_273601 & E_273833) ;
  assign /* unsigned    bit */  E_273877 = (E_273604 & E_273834) ;
  assign /* unsigned    bit */  E_273876 = (E_273588 & E_273751) ;
  assign /* unsigned    bit */  E_273875 = (E_273592 & E_273752) ;
  assign /* unsigned    bit */  E_273874 = (E_273595 & E_273753) ;
  assign /* unsigned    bit */  E_273873 = (E_273598 & E_273754) ;
  assign /* unsigned    bit */  E_273872 = (E_273601 & E_273755) ;
  assign /* unsigned    bit */  E_273871 = (E_273604 & E_273756) ;
  assign /* unsigned    bit */  E_273870 = (E_273588 & E_273808) ;
  assign /* unsigned    bit */  E_273869 = (E_273592 & E_273809) ;
  assign /* unsigned    bit */  E_273868 = (E_273595 & E_273810) ;
  assign /* unsigned    bit */  E_273867 = (E_273598 & E_273811) ;
  assign /* unsigned    bit */  E_273866 = (E_273601 & E_273812) ;
  assign /* unsigned    bit */  E_273865 = (E_273604 & E_273813) ;
  assign /* unsigned    bit */  E_273864 = (E_273588 & E_273762) ;
  assign /* unsigned    bit */  E_273863 = (E_273592 & E_273763) ;
  assign /* unsigned    bit */  E_273862 = (E_273595 & E_273764) ;
  assign /* unsigned    bit */  E_273861 = (E_273598 & E_273765) ;
  assign /* unsigned    bit */  E_273860 = (E_273601 & E_273766) ;
  assign /* unsigned    bit */  E_273859 = (E_273604 & E_273767) ;
  assign /* unsigned    bit */  E_273858 = (E_273588 & E_273590) ;
  assign /* unsigned    bit */  E_273857 = (E_273592 & E_273593) ;
  assign /* unsigned    bit */  E_273856 = (E_273595 & E_273596) ;
  assign /* unsigned    bit */  E_273855 = (E_273598 & E_273599) ;
  assign /* unsigned    bit */  E_273854 = (E_273601 & E_273602) ;
  assign /* unsigned    bit */  E_273853 = (E_273604 & E_273605) ;
  assign /* unsigned    bit */  E_273852 = (E_273623 & E_273695) ;
  assign /* unsigned    bit */  E_273851 = (E_273583 & E_273738) ;
  assign /* unsigned    bit */  E_273850 = (E_273837 & E_273734) ;
  assign /* unsigned    bit */  E_273849 = (E_273736 & E_273737) ;
  assign /* unsigned    bit */  E_273848 = (E_273604 & E_273747) ;
  assign /* unsigned    bit */  E_273847 = (E_273583 & E_273795) ;
  assign /* unsigned    bit */  E_273846 = (E_273837 & E_273793) ;
  assign /* unsigned    bit */  E_273845 = (E_273736 & E_273794) ;
  assign /* unsigned    bit */  E_273844 = (E_273604 & E_273804) ;
  assign /* unsigned    bit */  E_273843 = (E_273583 & E_273772) ;
  assign /* unsigned    bit */  E_273842 = (E_273837 & E_273770) ;
  assign /* unsigned    bit */  E_273841 = (E_273736 & E_273771) ;
  assign /* unsigned    bit */  E_273840 = (E_273604 & E_273781) ;
  assign /* unsigned    bit */  E_273839 = (E_273583 & E_273827) ;
  assign /* unsigned    bit */  E_273838 = (E_273735 & E_273826) ;
  assign /* unsigned    bit */  E_273837 = ( !E_273733 ) ;
  assign /* unsigned    bit */  E_273836 = (E_273837 & E_273838) ;
  assign /* unsigned    bit */  E_273835 = (E_273603 & E_273824) ;
  assign /* unsigned    bit */  E_273834 = (E_273614 & E_273651) ;
  assign /* unsigned    bit */  E_273833 = (E_273603 & E_273834) ;
  assign /* unsigned    bit */  E_273832 = (E_273600 & E_273833) ;
  assign /* unsigned    bit */  E_273831 = (E_273597 & E_273832) ;
  assign /* unsigned    bit */  E_273830 = (E_273594 & E_273831) ;
  assign /* unsigned    bit */  E_273829 = (E_273591 & E_273830) ;
  assign /* unsigned    bit */  E_273828 = (E_273587 & E_273829) ;
  assign /* unsigned    bit */  E_273827 = (E_273828 | E_273835) ;
  assign /* unsigned    bit */  E_273826 = (E_273584 & E_273827) ;
  assign /* unsigned    bit */  E_273825 = (E_273736 & E_273826) ;
  assign /* unsigned    bit */  E_273824 = (E_273614 & E_273709) ;
  assign /* unsigned    bit */  E_273823 = (E_273604 & E_273824) ;
  assign /* unsigned    bit */  E_273822 = (E_273583 & E_273749) ;
  assign /* unsigned    bit */  E_273821 = (E_273816 & E_273728) ;
  assign /* unsigned    bit */  E_273820 = (E_273730 & E_273731) ;
  assign /* unsigned    bit */  E_273819 = (E_273604 & E_273758) ;
  assign /* unsigned    bit */  E_273818 = (E_273583 & E_273806) ;
  assign /* unsigned    bit */  E_273817 = (E_273729 & E_273791) ;
  assign /* unsigned    bit */  E_273816 = ( !E_273727 ) ;
  assign /* unsigned    bit */  E_273815 = (E_273816 & E_273817) ;
  assign /* unsigned    bit */  E_273814 = (E_273603 & E_273789) ;
  assign /* unsigned    bit */  E_273813 = (E_273614 & E_273645) ;
  assign /* unsigned    bit */  E_273812 = (E_273603 & E_273813) ;
  assign /* unsigned    bit */  E_273811 = (E_273600 & E_273812) ;
  assign /* unsigned    bit */  E_273810 = (E_273597 & E_273811) ;
  assign /* unsigned    bit */  E_273809 = (E_273594 & E_273810) ;
  assign /* unsigned    bit */  E_273808 = (E_273591 & E_273809) ;
  assign /* unsigned    bit */  E_273807 = (E_273587 & E_273808) ;
  assign /* unsigned    bit */  E_273806 = (E_273807 | E_273814) ;
  assign /* unsigned    bit */  E_273805 = (E_273584 & E_273806) ;
  assign /* unsigned    bit */  E_273804 = (E_273614 & E_273715) ;
  assign /* unsigned    bit */  E_273803 = (E_273603 & E_273804) ;
  assign /* unsigned    bit */  E_273802 = (E_273614 & E_273658) ;
  assign /* unsigned    bit */  E_273801 = (E_273603 & E_273802) ;
  assign /* unsigned    bit */  E_273800 = (E_273600 & E_273801) ;
  assign /* unsigned    bit */  E_273799 = (E_273597 & E_273800) ;
  assign /* unsigned    bit */  E_273798 = (E_273594 & E_273799) ;
  assign /* unsigned    bit */  E_273797 = (E_273591 & E_273798) ;
  assign /* unsigned    bit */  E_273796 = (E_273587 & E_273797) ;
  assign /* unsigned    bit */  E_273795 = (E_273796 | E_273803) ;
  assign /* unsigned    bit */  E_273794 = (E_273584 & E_273795) ;
  assign /* unsigned    bit */  E_273793 = (E_273735 & E_273794) ;
  assign /* unsigned    bit */  E_273792 = (E_273733 & E_273793) ;
  assign /* unsigned    bit */  E_273791 = (E_273792 | E_273805) ;
  assign /* unsigned    bit */  E_273790 = (E_273730 & E_273791) ;
  assign /* unsigned    bit */  E_273789 = (E_273614 & E_273704) ;
  assign /* unsigned    bit */  E_273788 = (E_273604 & E_273789) ;
  assign /* unsigned    bit */  E_273787 = (E_273583 & E_273760) ;
  assign /* unsigned    bit */  E_273786 = ( !E_273723 ) ;
  assign /* unsigned    bit */  E_273785 = (E_273786 & E_273724) ;
  assign /* unsigned    bit */  E_273783 = ( !E_273784 ) ;
  assign /* unsigned    bit */  E_273782 = (E_273783 & E_273785) ;
  assign /* unsigned    bit */  E_273781 = (E_273614 & E_273713) ;
  assign /* unsigned    bit */  E_273780 = (E_273603 & E_273781) ;
  assign /* unsigned    bit */  E_273779 = (E_273614 & E_273656) ;
  assign /* unsigned    bit */  E_273778 = (E_273603 & E_273779) ;
  assign /* unsigned    bit */  E_273777 = (E_273600 & E_273778) ;
  assign /* unsigned    bit */  E_273776 = (E_273597 & E_273777) ;
  assign /* unsigned    bit */  E_273775 = (E_273594 & E_273776) ;
  assign /* unsigned    bit */  E_273774 = (E_273591 & E_273775) ;
  assign /* unsigned    bit */  E_273773 = (E_273587 & E_273774) ;
  assign /* unsigned    bit */  E_273772 = (E_273773 | E_273780) ;
  assign /* unsigned    bit */  E_273771 = (E_273584 & E_273772) ;
  assign /* unsigned    bit */  E_273770 = (E_273735 & E_273771) ;
  assign /* unsigned    bit */  E_273769 = (E_273733 & E_273770) ;
  assign /* unsigned    bit */  E_273768 = (E_273603 & E_273721) ;
  assign /* unsigned    bit */  E_273767 = (E_273614 & E_273615) ;
  assign /* unsigned    bit */  E_273766 = (E_273603 & E_273767) ;
  assign /* unsigned    bit */  E_273765 = (E_273600 & E_273766) ;
  assign /* unsigned    bit */  E_273764 = (E_273597 & E_273765) ;
  assign /* unsigned    bit */  E_273763 = (E_273594 & E_273764) ;
  assign /* unsigned    bit */  E_273762 = (E_273591 & E_273763) ;
  assign /* unsigned    bit */  E_273761 = (E_273587 & E_273762) ;
  assign /* unsigned    bit */  E_273760 = (E_273761 | E_273768) ;
  assign /* unsigned    bit */  E_273759 = (E_273584 & E_273760) ;
  assign /* unsigned    bit */  E_273758 = (E_273614 & E_273707) ;
  assign /* unsigned    bit */  E_273757 = (E_273603 & E_273758) ;
  assign /* unsigned    bit */  E_273756 = (E_273614 & E_273649) ;
  assign /* unsigned    bit */  E_273755 = (E_273603 & E_273756) ;
  assign /* unsigned    bit */  E_273754 = (E_273600 & E_273755) ;
  assign /* unsigned    bit */  E_273753 = (E_273597 & E_273754) ;
  assign /* unsigned    bit */  E_273752 = (E_273594 & E_273753) ;
  assign /* unsigned    bit */  E_273751 = (E_273591 & E_273752) ;
  assign /* unsigned    bit */  E_273750 = (E_273587 & E_273751) ;
  assign /* unsigned    bit */  E_273749 = (E_273750 | E_273757) ;
  assign /* unsigned    bit */  E_273748 = (E_273584 & E_273749) ;
  assign /* unsigned    bit */  E_273747 = (E_273614 & E_273718) ;
  assign /* unsigned    bit */  E_273746 = (E_273603 & E_273747) ;
  assign /* unsigned    bit */  E_273745 = (E_273614 & E_273661) ;
  assign /* unsigned    bit */  E_273744 = (E_273603 & E_273745) ;
  assign /* unsigned    bit */  E_273743 = (E_273600 & E_273744) ;
  assign /* unsigned    bit */  E_273742 = (E_273597 & E_273743) ;
  assign /* unsigned    bit */  E_273741 = (E_273594 & E_273742) ;
  assign /* unsigned    bit */  E_273740 = (E_273591 & E_273741) ;
  assign /* unsigned    bit */  E_273739 = (E_273587 & E_273740) ;
  assign /* unsigned    bit */  E_273738 = (E_273739 | E_273746) ;
  assign /* unsigned    bit */  E_273737 = (E_273584 & E_273738) ;
  assign /* unsigned    bit */  E_273735 = ( !E_273736 ) ;
  assign /* unsigned    bit */  E_273734 = (E_273735 & E_273737) ;
  assign /* unsigned    bit */  E_273732 = (E_273733 & E_273734) ;
  assign /* unsigned    bit */  E_273731 = (E_273732 | E_273748) ;
  assign /* unsigned    bit */  E_273729 = ( !E_273730 ) ;
  assign /* unsigned    bit */  E_273728 = (E_273729 & E_273731) ;
  assign /* unsigned    bit */  E_273726 = (E_273727 & E_273728) ;
  assign /* unsigned    bit */  E_273725 = (E_273726 | E_273759) ;
  assign /* unsigned    bit */  E_273724 = (E_273725 | E_273769) ;
  assign /* unsigned    bit */  E_273722 = (E_273723 & E_273724) ;
  assign /* unsigned    bit */  E_273721 = (E_273614 & E_273671) ;
  assign /* unsigned    bit */  E_273720 = (E_273604 & E_273721) ;
  assign /* unsigned    bit */  E_273719 = (E_273604 & E_273663) ;
  assign /* unsigned    bit */  E_273718 = (E_273616 & E_273716) ;
  assign /* unsigned    bit */  E_273717 = (E_273613 & E_273718) ;
  assign /* unsigned    bit */  E_273716 = (E_273647 & E_273711) ;
  assign /* unsigned    bit */  E_273715 = (E_273617 & E_273716) ;
  assign /* unsigned    bit */  E_273714 = (E_273613 & E_273715) ;
  assign /* unsigned    bit */  E_273713 = (E_273616 & E_273710) ;
  assign /* unsigned    bit */  E_273712 = (E_273613 & E_273713) ;
  assign /* unsigned    bit */  E_273711 = (E_273654 & E_273674) ;
  assign /* unsigned    bit */  E_273710 = (E_273619 & E_273711) ;
  assign /* unsigned    bit */  E_273709 = (E_273617 & E_273710) ;
  assign /* unsigned    bit */  E_273708 = (E_273613 & E_273709) ;
  assign /* unsigned    bit */  E_273707 = (E_273616 & E_273705) ;
  assign /* unsigned    bit */  E_273706 = (E_273613 & E_273707) ;
  assign /* unsigned    bit */  E_273705 = (E_273647 & E_273673) ;
  assign /* unsigned    bit */  E_273704 = (E_273617 & E_273705) ;
  assign /* unsigned    bit */  E_273703 = (E_273613 & E_273704) ;
  assign /* unsigned    bit */  E_273702 = (E_273617 & E_273672) ;
  assign /* unsigned    bit */  E_273701 = (E_273624 & E_273625) ;
  assign /* unsigned    bit */  E_273700 = (E_273627 & E_273629) ;
  assign /* unsigned    bit */  E_273699 = (E_273631 & E_273632) ;
  assign /* unsigned    bit */  E_273698 = (E_273634 & E_273635) ;
  assign /* unsigned    bit */  E_273697 = (E_273637 & E_273638) ;
  assign /* unsigned    bit */  E_273696 = (E_273640 & E_273641) ;
  assign /* unsigned    bit */  E_273695 = (E_273626 & E_273693) ;
  assign /* unsigned    bit */  E_273694 = (E_273624 & E_273695) ;
  assign /* unsigned    bit */  E_273693 = (E_273630 & E_273691) ;
  assign /* unsigned    bit */  E_273692 = (E_273627 & E_273693) ;
  assign /* unsigned    bit */  E_273691 = (E_273633 & E_273689) ;
  assign /* unsigned    bit */  E_273690 = (E_273631 & E_273691) ;
  assign /* unsigned    bit */  E_273689 = (E_273636 & E_273686) ;
  assign /* unsigned    bit */  E_273688 = (E_273634 & E_273689) ;
  assign /* unsigned    bit */  E_273687 = (E_273640 & E_273642) ;
  assign /* unsigned    bit */  E_273686 = (E_273639 & E_273642) ;
  assign /* unsigned    bit */  E_273685 = (E_273637 & E_273686) ;
  assign /* unsigned    bit */  E_273684 = (E_273685 | E_273687) ;
  assign /* unsigned    bit */  E_273683 = (E_273684 | E_273688) ;
  assign /* unsigned    bit */  E_273682 = (E_273683 | E_273690) ;
  assign /* unsigned    bit */  E_273681 = (E_273682 | E_273692) ;
  assign /* unsigned    bit */  E_273680 = (E_273681 | E_273694) ;
  assign /* unsigned    bit */  E_273679 = (E_273680 | E_273696) ;
  assign /* unsigned    bit */  E_273678 = (E_273679 | E_273697) ;
  assign /* unsigned    bit */  E_273677 = (E_273678 | E_273698) ;
  assign /* unsigned    bit */  E_273676 = (E_273677 | E_273699) ;
  assign /* unsigned    bit */  E_273675 = (E_273676 | E_273700) ;
  assign /* unsigned    bit */  E_273674 = (E_273675 | E_273701) ;
  assign /* unsigned    bit */  E_273673 = (E_273621 & E_273674) ;
  assign /* unsigned    bit */  E_273672 = (E_273619 & E_273673) ;
  assign /* unsigned    bit */  E_273671 = (E_273616 & E_273672) ;
  assign /* unsigned    bit */  E_273670 = (E_273613 & E_273671) ;
  assign /* unsigned    bit */  E_273669 = (E_273670 | E_273702) ;
  assign /* unsigned    bit */  E_273668 = (E_273669 | E_273703) ;
  assign /* unsigned    bit */  E_273667 = (E_273668 | E_273706) ;
  assign /* unsigned    bit */  E_273666 = (E_273667 | E_273708) ;
  assign /* unsigned    bit */  E_273665 = (E_273666 | E_273712) ;
  assign /* unsigned    bit */  E_273664 = (E_273665 | E_273714) ;
  assign /* unsigned    bit */  E_273663 = (E_273664 | E_273717) ;
  assign /* unsigned    bit */  E_273662 = (E_273603 & E_273663) ;
  assign /* unsigned    bit */  E_273661 = (E_273616 & E_273659) ;
  assign /* unsigned    bit */  E_273660 = (E_273613 & E_273661) ;
  assign /* unsigned    bit */  E_273659 = (E_273647 & E_273653) ;
  assign /* unsigned    bit */  E_273658 = (E_273617 & E_273659) ;
  assign /* unsigned    bit */  E_273657 = (E_273613 & E_273658) ;
  assign /* unsigned    bit */  E_273656 = (E_273616 & E_273652) ;
  assign /* unsigned    bit */  E_273655 = (E_273613 & E_273656) ;
  assign /* unsigned    bit */  E_273654 = ( !E_273621 ) ;
  assign /* unsigned    bit */  E_273653 = (E_273654 & E_273622) ;
  assign /* unsigned    bit */  E_273652 = (E_273619 & E_273653) ;
  assign /* unsigned    bit */  E_273651 = (E_273617 & E_273652) ;
  assign /* unsigned    bit */  E_273650 = (E_273613 & E_273651) ;
  assign /* unsigned    bit */  E_273649 = (E_273616 & E_273646) ;
  assign /* unsigned    bit */  E_273648 = (E_273613 & E_273649) ;
  assign /* unsigned    bit */  E_273647 = ( !E_273619 ) ;
  assign /* unsigned    bit */  E_273646 = (E_273647 & E_273620) ;
  assign /* unsigned    bit */  E_273645 = (E_273617 & E_273646) ;
  assign /* unsigned    bit */  E_273644 = (E_273613 & E_273645) ;
  assign /* unsigned    bit */  E_273643 = (E_273617 & E_273618) ;
  assign /* unsigned    bit */  E_273641 = ( !E_273642 ) ;
  assign /* unsigned    bit */  E_273640 = E_273628 [2]  ;
  assign /* unsigned    bit */  E_273639 = ( !E_273640 ) ;
  assign /* unsigned    bit */  E_273638 = (E_273639 & E_273641) ;
  assign /* unsigned    bit */  E_273637 = E_273628 [1]  ;
  assign /* unsigned    bit */  E_273636 = ( !E_273637 ) ;
  assign /* unsigned    bit */  E_273635 = (E_273636 & E_273638) ;
  assign /* unsigned    bit */  E_273634 = E_273628 [0]  ;
  assign /* unsigned    bit */  E_273633 = ( !E_273634 ) ;
  assign /* unsigned    bit */  E_273632 = (E_273633 & E_273635) ;
  assign /* unsigned    bit */  E_273631 = E_273628 [3]  ;
  assign /* unsigned    bit */  E_273630 = ( !E_273631 ) ;
  assign /* unsigned    bit */  E_273629 = (E_273630 & E_273632) ;
  assign /* unsigned    bit */  E_273627 = E_273628 [4]  ;
  assign /* unsigned    bit */  E_273626 = ( !E_273627 ) ;
  assign /* unsigned    bit */  E_273625 = (E_273626 & E_273629) ;
  assign /* unsigned    bit */  E_273623 = ( !E_273624 ) ;
  assign /* unsigned    bit */  E_273622 = (E_273623 & E_273625) ;
  assign /* unsigned    bit */  E_273620 = (E_273621 & E_273622) ;
  assign /* unsigned    bit */  E_273618 = (E_273619 & E_273620) ;
  assign /* unsigned    bit */  E_273616 = ( !E_273617 ) ;
  assign /* unsigned    bit */  E_273615 = (E_273616 & E_273618) ;
  assign /* unsigned    bit */  E_273613 = ( !E_273614 ) ;
  assign /* unsigned    bit */  E_273612 = (E_273613 & E_273615) ;
  assign /* unsigned    bit */  E_273611 = (E_273612 | E_273643) ;
  assign /* unsigned    bit */  E_273610 = (E_273611 | E_273644) ;
  assign /* unsigned    bit */  E_273609 = (E_273610 | E_273648) ;
  assign /* unsigned    bit */  E_273608 = (E_273609 | E_273650) ;
  assign /* unsigned    bit */  E_273607 = (E_273608 | E_273655) ;
  assign /* unsigned    bit */  E_273606 = (E_273607 | E_273657) ;
  assign /* unsigned    bit */  E_273605 = (E_273606 | E_273660) ;
  assign /* unsigned    bit */  E_273603 = ( !E_273604 ) ;
  assign /* unsigned    bit */  E_273602 = (E_273603 & E_273605) ;
  assign /* unsigned    bit */  E_273601 = E_273589 [4]  ;
  assign /* unsigned    bit */  E_273600 = ( !E_273601 ) ;
  assign /* unsigned    bit */  E_273599 = (E_273600 & E_273602) ;
  assign /* unsigned    bit */  E_273598 = E_273589 [3]  ;
  assign /* unsigned    bit */  E_273597 = ( !E_273598 ) ;
  assign /* unsigned    bit */  E_273596 = (E_273597 & E_273599) ;
  assign /* unsigned    bit */  E_273595 = E_273589 [0]  ;
  assign /* unsigned    bit */  E_273594 = ( !E_273595 ) ;
  assign /* unsigned    bit */  E_273593 = (E_273594 & E_273596) ;
  assign /* unsigned    bit */  E_273592 = E_273589 [1]  ;
  assign /* unsigned    bit */  E_273591 = ( !E_273592 ) ;
  assign /* unsigned    bit */  E_273590 = (E_273591 & E_273593) ;
  assign /* unsigned    bit */  E_273588 = E_273589 [2]  ;
  assign /* unsigned    bit */  E_273587 = ( !E_273588 ) ;
  assign /* unsigned    bit */  E_273586 = (E_273587 & E_273590) ;
  assign /* unsigned    bit */  E_273585 = (E_273586 | E_273662) ;
  assign /* unsigned    bit */  E_273583 = ( ~E_273584 ) ;
  assign /* unsigned    bit */  E_273582 = (E_273583 & E_273585) ;
  assign /* unsigned    bit */  E_273581 = (E_273582 | E_273719) ;
  assign /* unsigned    bit */  E_273580 = (E_273581 | E_273720) ;
  assign /* unsigned    bit */  E_273579 = (E_273580 | E_273722) ;
  assign /* unsigned    bit */  E_273578 = (E_273579 | E_273782) ;
  assign /* unsigned    bit */  E_273577 = (E_273578 | E_273787) ;
  assign /* unsigned    bit */  E_273576 = (E_273577 | E_273788) ;
  assign /* unsigned    bit */  E_273575 = (E_273576 | E_273790) ;
  assign /* unsigned    bit */  E_273574 = (E_273575 | E_273815) ;
  assign /* unsigned    bit */  E_273573 = (E_273574 | E_273818) ;
  assign /* unsigned    bit */  E_273572 = (E_273573 | E_273819) ;
  assign /* unsigned    bit */  E_273571 = (E_273572 | E_273820) ;
  assign /* unsigned    bit */  E_273570 = (E_273571 | E_273821) ;
  assign /* unsigned    bit */  E_273569 = (E_273570 | E_273822) ;
  assign /* unsigned    bit */  E_273568 = (E_273569 | E_273823) ;
  assign /* unsigned    bit */  E_273567 = (E_273568 | E_273825) ;
  assign /* unsigned    bit */  E_273566 = (E_273567 | E_273836) ;
  assign /* unsigned    bit */  E_273565 = (E_273566 | E_273839) ;
  assign /* unsigned    bit */  E_273564 = (E_273565 | E_273840) ;
  assign /* unsigned    bit */  E_273563 = (E_273564 | E_273841) ;
  assign /* unsigned    bit */  E_273562 = (E_273563 | E_273842) ;
  assign /* unsigned    bit */  E_273561 = (E_273562 | E_273843) ;
  assign /* unsigned    bit */  E_273560 = (E_273561 | E_273844) ;
  assign /* unsigned    bit */  E_273559 = (E_273560 | E_273845) ;
  assign /* unsigned    bit */  E_273558 = (E_273559 | E_273846) ;
  assign /* unsigned    bit */  E_273557 = (E_273558 | E_273847) ;
  assign /* unsigned    bit */  E_273556 = (E_273557 | E_273848) ;
  assign /* unsigned    bit */  E_273555 = (E_273556 | E_273849) ;
  assign /* unsigned    bit */  E_273554 = (E_273555 | E_273850) ;
  assign /* unsigned    bit */  E_273553 = (E_273554 | E_273851) ;
  assign /* unsigned    bit */  E_273552 = (E_273553 | E_273852) ;
  assign /* unsigned    bit */  E_273551 = (E_273552 | E_273853) ;
  assign /* unsigned    bit */  E_273550 = (E_273551 | E_273854) ;
  assign /* unsigned    bit */  E_273549 = (E_273550 | E_273855) ;
  assign /* unsigned    bit */  E_273548 = (E_273549 | E_273856) ;
  assign /* unsigned    bit */  E_273547 = (E_273548 | E_273857) ;
  assign /* unsigned    bit */  E_273546 = (E_273547 | E_273858) ;
  assign /* unsigned    bit */  E_273545 = (E_273546 | E_273859) ;
  assign /* unsigned    bit */  E_273544 = (E_273545 | E_273860) ;
  assign /* unsigned    bit */  E_273543 = (E_273544 | E_273861) ;
  assign /* unsigned    bit */  E_273542 = (E_273543 | E_273862) ;
  assign /* unsigned    bit */  E_273541 = (E_273542 | E_273863) ;
  assign /* unsigned    bit */  E_273540 = (E_273541 | E_273864) ;
  assign /* unsigned    bit */  E_273539 = (E_273540 | E_273865) ;
  assign /* unsigned    bit */  E_273538 = (E_273539 | E_273866) ;
  assign /* unsigned    bit */  E_273537 = (E_273538 | E_273867) ;
  assign /* unsigned    bit */  E_273536 = (E_273537 | E_273868) ;
  assign /* unsigned    bit */  E_273535 = (E_273536 | E_273869) ;
  assign /* unsigned    bit */  E_273534 = (E_273535 | E_273870) ;
  assign /* unsigned    bit */  E_273533 = (E_273534 | E_273871) ;
  assign /* unsigned    bit */  E_273532 = (E_273533 | E_273872) ;
  assign /* unsigned    bit */  E_273531 = (E_273532 | E_273873) ;
  assign /* unsigned    bit */  E_273530 = (E_273531 | E_273874) ;
  assign /* unsigned    bit */  E_273529 = (E_273530 | E_273875) ;
  assign /* unsigned    bit */  E_273528 = (E_273529 | E_273876) ;
  assign /* unsigned    bit */  E_273527 = (E_273528 | E_273877) ;
  assign /* unsigned    bit */  E_273526 = (E_273527 | E_273878) ;
  assign /* unsigned    bit */  E_273525 = (E_273526 | E_273879) ;
  assign /* unsigned    bit */  E_273524 = (E_273525 | E_273880) ;
  assign /* unsigned    bit */  E_273523 = (E_273524 | E_273881) ;
  assign /* unsigned    bit */  E_273522 = (E_273523 | E_273882) ;
  assign /* unsigned    bit */  E_273521 = (E_273522 | E_273883) ;
  assign /* unsigned    bit */  E_273520 = (E_273521 | E_273884) ;
  assign /* unsigned    bit */  E_273519 = (E_273520 | E_273885) ;
  assign /* unsigned    bit */  E_273518 = (E_273519 | E_273886) ;
  assign /* unsigned    bit */  E_273517 = (E_273518 | E_273887) ;
  assign /* unsigned    bit */  E_273516 = (E_273517 | E_273888) ;
  assign /* unsigned    bit */  E_273515 = (E_273516 | E_273889) ;
  assign /* unsigned    bit */  E_273514 = (E_273515 | E_273890) ;
  assign /* unsigned    bit */  E_273513 = (E_273514 | E_273891) ;
  assign /* unsigned    bit */  E_273512 = (E_273513 | E_273892) ;
  assign /* unsigned    bit */  E_273511 = (E_273512 | E_273893) ;
  assign /* unsigned    bit */  E_273510 = (E_273511 | E_273894) ;
  assign /* unsigned    bit */  E_273509 = (E_273510 | E_273895) ;
  assign /* unsigned    bit */  E_273508 = (E_273509 | E_273896) ;
  assign /* unsigned    bit */  E_273507 = (E_273508 | E_273897) ;
  assign /* unsigned    bit */  E_273506 = (E_273507 | E_273898) ;
  assign /* unsigned    bit */  E_273505 = (E_273506 | E_273899) ;
  assign /* unsigned    bit */  E_273504 = (E_273505 | E_273900) ;
  assign /* unsigned    bit */  E_273502 = ( !E_273503 ) ;
  assign /* unsigned    bit */  E_273501 = (E_273502 & E_273504) ;
  assign /* unsigned    bit */  E_273499 = (E_273500 & E_273501) ;
  assign /* unsigned    bit */  E_273497 = ( !E_273498 ) ;
  assign /* unsigned    bit */  E_273496 = (E_273497 | E_273499) ;
endmodule



//Hier for 'O_write_data_data_sva'
module temp_odc_impl_1452 ( reg_W_instr_in_rsci_oswt_cse_1_0 , land_9_lpi_1_dfm_1_1_1
 , t_out ) ;
 input wire  reg_W_instr_in_rsci_oswt_cse_1_0 ; 
 input wire  land_9_lpi_1_dfm_1_1_1 ; 
 output wire  t_out ; 
 wire E_273906 ; 
assign t_out = E_273906 ;
 wire E_273905 ; 
assign E_273905 = land_9_lpi_1_dfm_1_1_1 ;
 wire E_273904 ; 
assign E_273904 = reg_W_instr_in_rsci_oswt_cse_1_0 ;
 wire E_273903 ; 
 wire E_273902 ; 
  assign /* unsigned    bit */  E_273906 = ( !E_273902 ) ;
  assign /* unsigned    bit */  E_273903 = ( !E_273904 ) ;
  assign /* unsigned    bit */  E_273902 = (E_273903 & E_273905) ;
endmodule



//Hier for 'O_wr_data_rsci_ivld_bfwt'
module temp_odc_impl_1453 ( O_wr_data_rsci_bcwt_0 , run_wten_1 , reg_O_wr_data_rsci_irdy_run_psct_cse_2
 , t_out ) ;
 input wire  O_wr_data_rsci_bcwt_0 ; 
 input wire  run_wten_1 ; 
 input wire  reg_O_wr_data_rsci_irdy_run_psct_cse_2 ; 
 output wire  t_out ; 
 wire E_273916 ; 
assign t_out = E_273916 ;
 wire E_273915 ; 
assign E_273915 = reg_O_wr_data_rsci_irdy_run_psct_cse_2 ;
 wire E_273914 ; 
 wire E_273913 ; 
assign E_273913 = run_wten_1 ;
 wire E_273912 ; 
 wire E_273911 ; 
 wire E_273910 ; 
 wire E_273909 ; 
assign E_273909 = O_wr_data_rsci_bcwt_0 ;
 wire E_273908 ; 
 wire E_273907 ; 
  assign /* unsigned    bit */  E_273916 = ( !E_273907 ) ;
  assign /* unsigned    bit */  E_273914 = ( !E_273915 ) ;
  assign /* unsigned    bit */  E_273912 = (E_273913 | E_273914) ;
  assign /* unsigned    bit */  E_273911 = (E_273909 | E_273912) ;
  assign /* unsigned    bit */  E_273910 = ( !E_273911 ) ;
  assign /* unsigned    bit */  E_273908 = ( ~E_273909 ) ;
  assign /* unsigned    bit */  E_273907 = (E_273908 | E_273910) ;
endmodule



//Hier for 'O_wr_data_rsci_idat_bfwt'
module temp_odc_impl_1454 ( O_wr_data_rsci_bcwt_0 , run_wten_1 , reg_O_wr_data_rsci_irdy_run_psct_cse_2
 , t_out ) ;
 input wire  O_wr_data_rsci_bcwt_0 ; 
 input wire  run_wten_1 ; 
 input wire  reg_O_wr_data_rsci_irdy_run_psct_cse_2 ; 
 output wire  t_out ; 
 wire E_273924 ; 
assign t_out = E_273924 ;
 wire E_273923 ; 
assign E_273923 = reg_O_wr_data_rsci_irdy_run_psct_cse_2 ;
 wire E_273922 ; 
 wire E_273921 ; 
assign E_273921 = run_wten_1 ;
 wire E_273920 ; 
 wire E_273919 ; 
assign E_273919 = O_wr_data_rsci_bcwt_0 ;
 wire E_273918 ; 
 wire E_273917 ; 
  assign /* unsigned    bit */  E_273924 = ( !E_273917 ) ;
  assign /* unsigned    bit */  E_273922 = ( !E_273923 ) ;
  assign /* unsigned    bit */  E_273920 = (E_273921 | E_273922) ;
  assign /* unsigned    bit */  E_273918 = (E_273919 | E_273920) ;
  assign /* unsigned    bit */  E_273917 = ( !E_273918 ) ;
endmodule



