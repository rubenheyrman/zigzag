VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO SRAM_128x1296_2P
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 536.256 BY 161.728 ;
  SYMMETRY X Y R90 ;

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 519.840 0.000 519.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 519.840 0.000 519.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 519.840 0.000 519.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 519.840 0.000 519.992 0.152 ;
    END
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 513.456 0.000 513.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 513.456 0.000 513.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 513.456 0.000 513.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 513.456 0.000 513.608 0.152 ;
    END
  END CSB1

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 507.072 0.000 507.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 507.072 0.000 507.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 507.072 0.000 507.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 507.072 0.000 507.224 0.152 ;
    END
  END OEB1

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 500.688 0.000 500.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 500.688 0.000 500.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 500.688 0.000 500.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 500.688 0.000 500.840 0.152 ;
    END
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 500.384 0.000 500.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 500.384 0.000 500.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 500.384 0.000 500.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 500.384 0.000 500.536 0.152 ;
    END
  END O1[2]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 500.080 0.000 500.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 500.080 0.000 500.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 500.080 0.000 500.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 500.080 0.000 500.232 0.152 ;
    END
  END O1[1]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 499.776 0.000 499.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 499.776 0.000 499.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 499.776 0.000 499.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 499.776 0.000 499.928 0.152 ;
    END
  END O1[0]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 493.392 0.000 493.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 493.392 0.000 493.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 493.392 0.000 493.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 493.392 0.000 493.544 0.152 ;
    END
  END O1[7]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 493.088 0.000 493.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 493.088 0.000 493.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 493.088 0.000 493.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 493.088 0.000 493.240 0.152 ;
    END
  END O1[6]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 492.784 0.000 492.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 492.784 0.000 492.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 492.784 0.000 492.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 492.784 0.000 492.936 0.152 ;
    END
  END O1[5]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 492.480 0.000 492.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 492.480 0.000 492.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 492.480 0.000 492.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 492.480 0.000 492.632 0.152 ;
    END
  END O1[4]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 486.096 0.000 486.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 486.096 0.000 486.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 486.096 0.000 486.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 486.096 0.000 486.248 0.152 ;
    END
  END O1[11]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 485.792 0.000 485.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 485.792 0.000 485.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 485.792 0.000 485.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 485.792 0.000 485.944 0.152 ;
    END
  END O1[10]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 485.488 0.000 485.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 485.488 0.000 485.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 485.488 0.000 485.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 485.488 0.000 485.640 0.152 ;
    END
  END O1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 485.184 0.000 485.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 485.184 0.000 485.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 485.184 0.000 485.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 485.184 0.000 485.336 0.152 ;
    END
  END O1[8]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 478.800 0.000 478.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 478.800 0.000 478.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 478.800 0.000 478.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 478.800 0.000 478.952 0.152 ;
    END
  END O1[15]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 478.496 0.000 478.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 478.496 0.000 478.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 478.496 0.000 478.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 478.496 0.000 478.648 0.152 ;
    END
  END O1[14]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 478.192 0.000 478.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 478.192 0.000 478.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 478.192 0.000 478.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 478.192 0.000 478.344 0.152 ;
    END
  END O1[13]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 477.888 0.000 478.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 477.888 0.000 478.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 477.888 0.000 478.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 477.888 0.000 478.040 0.152 ;
    END
  END O1[12]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 471.504 0.000 471.656 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 471.504 0.000 471.656 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 471.504 0.000 471.656 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 471.504 0.000 471.656 0.152 ;
    END
  END O1[19]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 471.200 0.000 471.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 471.200 0.000 471.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 471.200 0.000 471.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 471.200 0.000 471.352 0.152 ;
    END
  END O1[18]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 470.896 0.000 471.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 470.896 0.000 471.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 470.896 0.000 471.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 470.896 0.000 471.048 0.152 ;
    END
  END O1[17]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 470.592 0.000 470.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 470.592 0.000 470.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 470.592 0.000 470.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 470.592 0.000 470.744 0.152 ;
    END
  END O1[16]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 464.208 0.000 464.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 464.208 0.000 464.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 464.208 0.000 464.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 464.208 0.000 464.360 0.152 ;
    END
  END O1[23]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 463.904 0.000 464.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 463.904 0.000 464.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 463.904 0.000 464.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 463.904 0.000 464.056 0.152 ;
    END
  END O1[22]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 463.600 0.000 463.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 463.600 0.000 463.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 463.600 0.000 463.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 463.600 0.000 463.752 0.152 ;
    END
  END O1[21]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 463.296 0.000 463.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 463.296 0.000 463.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 463.296 0.000 463.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 463.296 0.000 463.448 0.152 ;
    END
  END O1[20]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 456.912 0.000 457.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 456.912 0.000 457.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 456.912 0.000 457.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 456.912 0.000 457.064 0.152 ;
    END
  END O1[27]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 456.608 0.000 456.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 456.608 0.000 456.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 456.608 0.000 456.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 456.608 0.000 456.760 0.152 ;
    END
  END O1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 456.304 0.000 456.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 456.304 0.000 456.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 456.304 0.000 456.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 456.304 0.000 456.456 0.152 ;
    END
  END O1[25]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 456.000 0.000 456.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 456.000 0.000 456.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 456.000 0.000 456.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 456.000 0.000 456.152 0.152 ;
    END
  END O1[24]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 449.616 0.000 449.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 449.616 0.000 449.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 449.616 0.000 449.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 449.616 0.000 449.768 0.152 ;
    END
  END O1[31]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 449.312 0.000 449.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 449.312 0.000 449.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 449.312 0.000 449.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 449.312 0.000 449.464 0.152 ;
    END
  END O1[30]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 449.008 0.000 449.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 449.008 0.000 449.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 449.008 0.000 449.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 449.008 0.000 449.160 0.152 ;
    END
  END O1[29]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 448.704 0.000 448.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 448.704 0.000 448.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 448.704 0.000 448.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 448.704 0.000 448.856 0.152 ;
    END
  END O1[28]

  PIN O1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 442.320 0.000 442.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 442.320 0.000 442.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 442.320 0.000 442.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 442.320 0.000 442.472 0.152 ;
    END
  END O1[35]

  PIN O1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 442.016 0.000 442.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 442.016 0.000 442.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 442.016 0.000 442.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 442.016 0.000 442.168 0.152 ;
    END
  END O1[34]

  PIN O1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 441.712 0.000 441.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 441.712 0.000 441.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 441.712 0.000 441.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 441.712 0.000 441.864 0.152 ;
    END
  END O1[33]

  PIN O1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 441.408 0.000 441.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 441.408 0.000 441.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 441.408 0.000 441.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 441.408 0.000 441.560 0.152 ;
    END
  END O1[32]

  PIN O1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.024 0.000 435.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 435.024 0.000 435.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 435.024 0.000 435.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 435.024 0.000 435.176 0.152 ;
    END
  END O1[39]

  PIN O1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 434.720 0.000 434.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 434.720 0.000 434.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 434.720 0.000 434.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 434.720 0.000 434.872 0.152 ;
    END
  END O1[38]

  PIN O1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 434.416 0.000 434.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 434.416 0.000 434.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 434.416 0.000 434.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 434.416 0.000 434.568 0.152 ;
    END
  END O1[37]

  PIN O1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 434.112 0.000 434.264 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 434.112 0.000 434.264 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 434.112 0.000 434.264 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 434.112 0.000 434.264 0.152 ;
    END
  END O1[36]

  PIN O1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.728 0.000 427.880 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 427.728 0.000 427.880 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 427.728 0.000 427.880 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 427.728 0.000 427.880 0.152 ;
    END
  END O1[43]

  PIN O1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.424 0.000 427.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 427.424 0.000 427.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 427.424 0.000 427.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 427.424 0.000 427.576 0.152 ;
    END
  END O1[42]

  PIN O1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.120 0.000 427.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 427.120 0.000 427.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 427.120 0.000 427.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 427.120 0.000 427.272 0.152 ;
    END
  END O1[41]

  PIN O1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 426.816 0.000 426.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 426.816 0.000 426.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 426.816 0.000 426.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 426.816 0.000 426.968 0.152 ;
    END
  END O1[40]

  PIN O1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.432 0.000 420.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 420.432 0.000 420.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 420.432 0.000 420.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 420.432 0.000 420.584 0.152 ;
    END
  END O1[47]

  PIN O1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.128 0.000 420.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 420.128 0.000 420.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 420.128 0.000 420.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 420.128 0.000 420.280 0.152 ;
    END
  END O1[46]

  PIN O1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 419.824 0.000 419.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 419.824 0.000 419.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 419.824 0.000 419.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 419.824 0.000 419.976 0.152 ;
    END
  END O1[45]

  PIN O1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 419.520 0.000 419.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 419.520 0.000 419.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 419.520 0.000 419.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 419.520 0.000 419.672 0.152 ;
    END
  END O1[44]

  PIN O1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 413.136 0.000 413.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 413.136 0.000 413.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 413.136 0.000 413.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 413.136 0.000 413.288 0.152 ;
    END
  END O1[51]

  PIN O1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.832 0.000 412.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 412.832 0.000 412.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 412.832 0.000 412.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 412.832 0.000 412.984 0.152 ;
    END
  END O1[50]

  PIN O1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.528 0.000 412.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 412.528 0.000 412.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 412.528 0.000 412.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 412.528 0.000 412.680 0.152 ;
    END
  END O1[49]

  PIN O1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.224 0.000 412.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 412.224 0.000 412.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 412.224 0.000 412.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 412.224 0.000 412.376 0.152 ;
    END
  END O1[48]

  PIN O1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 405.840 0.000 405.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 405.840 0.000 405.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 405.840 0.000 405.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 405.840 0.000 405.992 0.152 ;
    END
  END O1[55]

  PIN O1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 405.536 0.000 405.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 405.536 0.000 405.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 405.536 0.000 405.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 405.536 0.000 405.688 0.152 ;
    END
  END O1[54]

  PIN O1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 405.232 0.000 405.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 405.232 0.000 405.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 405.232 0.000 405.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 405.232 0.000 405.384 0.152 ;
    END
  END O1[53]

  PIN O1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 404.928 0.000 405.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 404.928 0.000 405.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 404.928 0.000 405.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 404.928 0.000 405.080 0.152 ;
    END
  END O1[52]

  PIN O1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 398.544 0.000 398.696 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 398.544 0.000 398.696 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 398.544 0.000 398.696 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 398.544 0.000 398.696 0.152 ;
    END
  END O1[59]

  PIN O1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 398.240 0.000 398.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 398.240 0.000 398.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 398.240 0.000 398.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 398.240 0.000 398.392 0.152 ;
    END
  END O1[58]

  PIN O1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 397.936 0.000 398.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 397.936 0.000 398.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 397.936 0.000 398.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 397.936 0.000 398.088 0.152 ;
    END
  END O1[57]

  PIN O1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 397.632 0.000 397.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 397.632 0.000 397.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 397.632 0.000 397.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 397.632 0.000 397.784 0.152 ;
    END
  END O1[56]

  PIN O1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 391.248 0.000 391.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 391.248 0.000 391.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 391.248 0.000 391.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 391.248 0.000 391.400 0.152 ;
    END
  END O1[63]

  PIN O1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.944 0.000 391.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 390.944 0.000 391.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 390.944 0.000 391.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 390.944 0.000 391.096 0.152 ;
    END
  END O1[62]

  PIN O1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.640 0.000 390.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 390.640 0.000 390.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 390.640 0.000 390.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 390.640 0.000 390.792 0.152 ;
    END
  END O1[61]

  PIN O1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.336 0.000 390.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 390.336 0.000 390.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 390.336 0.000 390.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 390.336 0.000 390.488 0.152 ;
    END
  END O1[60]

  PIN O1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.952 0.000 384.104 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 383.952 0.000 384.104 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 383.952 0.000 384.104 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 383.952 0.000 384.104 0.152 ;
    END
  END O1[67]

  PIN O1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.648 0.000 383.800 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 383.648 0.000 383.800 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 383.648 0.000 383.800 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 383.648 0.000 383.800 0.152 ;
    END
  END O1[66]

  PIN O1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.344 0.000 383.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 383.344 0.000 383.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 383.344 0.000 383.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 383.344 0.000 383.496 0.152 ;
    END
  END O1[65]

  PIN O1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.040 0.000 383.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 383.040 0.000 383.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 383.040 0.000 383.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 383.040 0.000 383.192 0.152 ;
    END
  END O1[64]

  PIN O1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.656 0.000 376.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 376.656 0.000 376.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 376.656 0.000 376.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 376.656 0.000 376.808 0.152 ;
    END
  END O1[71]

  PIN O1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.352 0.000 376.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 376.352 0.000 376.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 376.352 0.000 376.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 376.352 0.000 376.504 0.152 ;
    END
  END O1[70]

  PIN O1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.048 0.000 376.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 376.048 0.000 376.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 376.048 0.000 376.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 376.048 0.000 376.200 0.152 ;
    END
  END O1[69]

  PIN O1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 375.744 0.000 375.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 375.744 0.000 375.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 375.744 0.000 375.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 375.744 0.000 375.896 0.152 ;
    END
  END O1[68]

  PIN O1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 369.360 0.000 369.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 369.360 0.000 369.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 369.360 0.000 369.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 369.360 0.000 369.512 0.152 ;
    END
  END O1[75]

  PIN O1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 369.056 0.000 369.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 369.056 0.000 369.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 369.056 0.000 369.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 369.056 0.000 369.208 0.152 ;
    END
  END O1[74]

  PIN O1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 368.752 0.000 368.904 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 368.752 0.000 368.904 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 368.752 0.000 368.904 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 368.752 0.000 368.904 0.152 ;
    END
  END O1[73]

  PIN O1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 368.448 0.000 368.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 368.448 0.000 368.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 368.448 0.000 368.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 368.448 0.000 368.600 0.152 ;
    END
  END O1[72]

  PIN O1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 362.064 0.000 362.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 362.064 0.000 362.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 362.064 0.000 362.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 362.064 0.000 362.216 0.152 ;
    END
  END O1[79]

  PIN O1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 361.760 0.000 361.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 361.760 0.000 361.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 361.760 0.000 361.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 361.760 0.000 361.912 0.152 ;
    END
  END O1[78]

  PIN O1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 361.456 0.000 361.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 361.456 0.000 361.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 361.456 0.000 361.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 361.456 0.000 361.608 0.152 ;
    END
  END O1[77]

  PIN O1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 361.152 0.000 361.304 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 361.152 0.000 361.304 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 361.152 0.000 361.304 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 361.152 0.000 361.304 0.152 ;
    END
  END O1[76]

  PIN O1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.768 0.000 354.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 354.768 0.000 354.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 354.768 0.000 354.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 354.768 0.000 354.920 0.152 ;
    END
  END O1[83]

  PIN O1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.464 0.000 354.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 354.464 0.000 354.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 354.464 0.000 354.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 354.464 0.000 354.616 0.152 ;
    END
  END O1[82]

  PIN O1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.160 0.000 354.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 354.160 0.000 354.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 354.160 0.000 354.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 354.160 0.000 354.312 0.152 ;
    END
  END O1[81]

  PIN O1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 353.856 0.000 354.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 353.856 0.000 354.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 353.856 0.000 354.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 353.856 0.000 354.008 0.152 ;
    END
  END O1[80]

  PIN O1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.472 0.000 347.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 347.472 0.000 347.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 347.472 0.000 347.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 347.472 0.000 347.624 0.152 ;
    END
  END O1[87]

  PIN O1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.168 0.000 347.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 347.168 0.000 347.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 347.168 0.000 347.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 347.168 0.000 347.320 0.152 ;
    END
  END O1[86]

  PIN O1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.864 0.000 347.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 346.864 0.000 347.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 346.864 0.000 347.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 346.864 0.000 347.016 0.152 ;
    END
  END O1[85]

  PIN O1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.560 0.000 346.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 346.560 0.000 346.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 346.560 0.000 346.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 346.560 0.000 346.712 0.152 ;
    END
  END O1[84]

  PIN O1[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.176 0.000 340.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 340.176 0.000 340.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 340.176 0.000 340.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 340.176 0.000 340.328 0.152 ;
    END
  END O1[91]

  PIN O1[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.872 0.000 340.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 339.872 0.000 340.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 339.872 0.000 340.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 339.872 0.000 340.024 0.152 ;
    END
  END O1[90]

  PIN O1[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.568 0.000 339.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 339.568 0.000 339.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 339.568 0.000 339.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 339.568 0.000 339.720 0.152 ;
    END
  END O1[89]

  PIN O1[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.264 0.000 339.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 339.264 0.000 339.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 339.264 0.000 339.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 339.264 0.000 339.416 0.152 ;
    END
  END O1[88]

  PIN O1[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.880 0.000 333.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 332.880 0.000 333.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 332.880 0.000 333.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 332.880 0.000 333.032 0.152 ;
    END
  END O1[95]

  PIN O1[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.576 0.000 332.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 332.576 0.000 332.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 332.576 0.000 332.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 332.576 0.000 332.728 0.152 ;
    END
  END O1[94]

  PIN O1[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.272 0.000 332.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 332.272 0.000 332.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 332.272 0.000 332.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 332.272 0.000 332.424 0.152 ;
    END
  END O1[93]

  PIN O1[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.968 0.000 332.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 331.968 0.000 332.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 331.968 0.000 332.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 331.968 0.000 332.120 0.152 ;
    END
  END O1[92]

  PIN O1[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.584 0.000 325.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 325.584 0.000 325.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 325.584 0.000 325.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 325.584 0.000 325.736 0.152 ;
    END
  END O1[99]

  PIN O1[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.280 0.000 325.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 325.280 0.000 325.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 325.280 0.000 325.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 325.280 0.000 325.432 0.152 ;
    END
  END O1[98]

  PIN O1[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.976 0.000 325.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 324.976 0.000 325.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 324.976 0.000 325.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 324.976 0.000 325.128 0.152 ;
    END
  END O1[97]

  PIN O1[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.672 0.000 324.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 324.672 0.000 324.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 324.672 0.000 324.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 324.672 0.000 324.824 0.152 ;
    END
  END O1[96]

  PIN O1[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.288 0.000 318.440 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 318.288 0.000 318.440 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 318.288 0.000 318.440 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 318.288 0.000 318.440 0.152 ;
    END
  END O1[103]

  PIN O1[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.984 0.000 318.136 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 317.984 0.000 318.136 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 317.984 0.000 318.136 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 317.984 0.000 318.136 0.152 ;
    END
  END O1[102]

  PIN O1[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.680 0.000 317.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 317.680 0.000 317.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 317.680 0.000 317.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 317.680 0.000 317.832 0.152 ;
    END
  END O1[101]

  PIN O1[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.376 0.000 317.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 317.376 0.000 317.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 317.376 0.000 317.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 317.376 0.000 317.528 0.152 ;
    END
  END O1[100]

  PIN O1[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.992 0.000 311.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 310.992 0.000 311.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 310.992 0.000 311.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 310.992 0.000 311.144 0.152 ;
    END
  END O1[107]

  PIN O1[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.688 0.000 310.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 310.688 0.000 310.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 310.688 0.000 310.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 310.688 0.000 310.840 0.152 ;
    END
  END O1[106]

  PIN O1[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.384 0.000 310.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 310.384 0.000 310.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 310.384 0.000 310.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 310.384 0.000 310.536 0.152 ;
    END
  END O1[105]

  PIN O1[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.080 0.000 310.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 310.080 0.000 310.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 310.080 0.000 310.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 310.080 0.000 310.232 0.152 ;
    END
  END O1[104]

  PIN O1[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.696 0.000 303.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 303.696 0.000 303.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 303.696 0.000 303.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 303.696 0.000 303.848 0.152 ;
    END
  END O1[111]

  PIN O1[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.392 0.000 303.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 303.392 0.000 303.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 303.392 0.000 303.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 303.392 0.000 303.544 0.152 ;
    END
  END O1[110]

  PIN O1[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.088 0.000 303.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 303.088 0.000 303.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 303.088 0.000 303.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 303.088 0.000 303.240 0.152 ;
    END
  END O1[109]

  PIN O1[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 302.784 0.000 302.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 302.784 0.000 302.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 302.784 0.000 302.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 302.784 0.000 302.936 0.152 ;
    END
  END O1[108]

  PIN O1[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 296.400 0.000 296.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 296.400 0.000 296.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 296.400 0.000 296.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 296.400 0.000 296.552 0.152 ;
    END
  END O1[115]

  PIN O1[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 296.096 0.000 296.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 296.096 0.000 296.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 296.096 0.000 296.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 296.096 0.000 296.248 0.152 ;
    END
  END O1[114]

  PIN O1[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.792 0.000 295.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 295.792 0.000 295.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 295.792 0.000 295.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 295.792 0.000 295.944 0.152 ;
    END
  END O1[113]

  PIN O1[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.488 0.000 295.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 295.488 0.000 295.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 295.488 0.000 295.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 295.488 0.000 295.640 0.152 ;
    END
  END O1[112]

  PIN O1[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 289.104 0.000 289.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 289.104 0.000 289.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 289.104 0.000 289.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 289.104 0.000 289.256 0.152 ;
    END
  END O1[119]

  PIN O1[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 288.800 0.000 288.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 288.800 0.000 288.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 288.800 0.000 288.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 288.800 0.000 288.952 0.152 ;
    END
  END O1[118]

  PIN O1[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 288.496 0.000 288.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 288.496 0.000 288.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 288.496 0.000 288.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 288.496 0.000 288.648 0.152 ;
    END
  END O1[117]

  PIN O1[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 288.192 0.000 288.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 288.192 0.000 288.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 288.192 0.000 288.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 288.192 0.000 288.344 0.152 ;
    END
  END O1[116]

  PIN O1[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 281.808 0.000 281.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 281.808 0.000 281.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 281.808 0.000 281.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 281.808 0.000 281.960 0.152 ;
    END
  END O1[123]

  PIN O1[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 281.504 0.000 281.656 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 281.504 0.000 281.656 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 281.504 0.000 281.656 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 281.504 0.000 281.656 0.152 ;
    END
  END O1[122]

  PIN O1[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 281.200 0.000 281.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 281.200 0.000 281.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 281.200 0.000 281.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 281.200 0.000 281.352 0.152 ;
    END
  END O1[121]

  PIN O1[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 280.896 0.000 281.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 280.896 0.000 281.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 280.896 0.000 281.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 280.896 0.000 281.048 0.152 ;
    END
  END O1[120]

  PIN O1[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 274.512 0.000 274.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 274.512 0.000 274.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 274.512 0.000 274.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 274.512 0.000 274.664 0.152 ;
    END
  END O1[127]

  PIN O1[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 274.208 0.000 274.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 274.208 0.000 274.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 274.208 0.000 274.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 274.208 0.000 274.360 0.152 ;
    END
  END O1[126]

  PIN O1[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 273.904 0.000 274.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 273.904 0.000 274.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 273.904 0.000 274.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 273.904 0.000 274.056 0.152 ;
    END
  END O1[125]

  PIN O1[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 273.600 0.000 273.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 273.600 0.000 273.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 273.600 0.000 273.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 273.600 0.000 273.752 0.152 ;
    END
  END O1[124]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.104 141.512 536.256 141.664 ;
    END
    PORT
      LAYER M3 ;
        RECT 536.104 141.512 536.256 141.664 ;
    END
    PORT
      LAYER M4 ;
        RECT 536.104 141.512 536.256 141.664 ;
    END
    PORT
      LAYER M5 ;
        RECT 536.104 141.512 536.256 141.664 ;
    END
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.104 137.864 536.256 138.016 ;
    END
    PORT
      LAYER M3 ;
        RECT 536.104 137.864 536.256 138.016 ;
    END
    PORT
      LAYER M4 ;
        RECT 536.104 137.864 536.256 138.016 ;
    END
    PORT
      LAYER M5 ;
        RECT 536.104 137.864 536.256 138.016 ;
    END
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.104 134.216 536.256 134.368 ;
    END
    PORT
      LAYER M3 ;
        RECT 536.104 134.216 536.256 134.368 ;
    END
    PORT
      LAYER M4 ;
        RECT 536.104 134.216 536.256 134.368 ;
    END
    PORT
      LAYER M5 ;
        RECT 536.104 134.216 536.256 134.368 ;
    END
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.104 130.568 536.256 130.720 ;
    END
    PORT
      LAYER M3 ;
        RECT 536.104 130.568 536.256 130.720 ;
    END
    PORT
      LAYER M4 ;
        RECT 536.104 130.568 536.256 130.720 ;
    END
    PORT
      LAYER M5 ;
        RECT 536.104 130.568 536.256 130.720 ;
    END
  END A1[3]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.104 126.920 536.256 127.072 ;
    END
    PORT
      LAYER M3 ;
        RECT 536.104 126.920 536.256 127.072 ;
    END
    PORT
      LAYER M4 ;
        RECT 536.104 126.920 536.256 127.072 ;
    END
    PORT
      LAYER M5 ;
        RECT 536.104 126.920 536.256 127.072 ;
    END
  END A1[4]

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.104 123.272 536.256 123.424 ;
    END
    PORT
      LAYER M3 ;
        RECT 536.104 123.272 536.256 123.424 ;
    END
    PORT
      LAYER M4 ;
        RECT 536.104 123.272 536.256 123.424 ;
    END
    PORT
      LAYER M5 ;
        RECT 536.104 123.272 536.256 123.424 ;
    END
  END A1[5]

  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.104 119.624 536.256 119.776 ;
    END
    PORT
      LAYER M3 ;
        RECT 536.104 119.624 536.256 119.776 ;
    END
    PORT
      LAYER M4 ;
        RECT 536.104 119.624 536.256 119.776 ;
    END
    PORT
      LAYER M5 ;
        RECT 536.104 119.624 536.256 119.776 ;
    END
  END A1[6]

  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.104 115.976 536.256 116.128 ;
    END
    PORT
      LAYER M3 ;
        RECT 536.104 115.976 536.256 116.128 ;
    END
    PORT
      LAYER M4 ;
        RECT 536.104 115.976 536.256 116.128 ;
    END
    PORT
      LAYER M5 ;
        RECT 536.104 115.976 536.256 116.128 ;
    END
  END A1[7]

  PIN A1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.104 112.328 536.256 112.480 ;
    END
    PORT
      LAYER M3 ;
        RECT 536.104 112.328 536.256 112.480 ;
    END
    PORT
      LAYER M4 ;
        RECT 536.104 112.328 536.256 112.480 ;
    END
    PORT
      LAYER M5 ;
        RECT 536.104 112.328 536.256 112.480 ;
    END
  END A1[8]

  PIN A1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.104 108.680 536.256 108.832 ;
    END
    PORT
      LAYER M3 ;
        RECT 536.104 108.680 536.256 108.832 ;
    END
    PORT
      LAYER M4 ;
        RECT 536.104 108.680 536.256 108.832 ;
    END
    PORT
      LAYER M5 ;
        RECT 536.104 108.680 536.256 108.832 ;
    END
  END A1[9]

  PIN A1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.104 105.032 536.256 105.184 ;
    END
    PORT
      LAYER M3 ;
        RECT 536.104 105.032 536.256 105.184 ;
    END
    PORT
      LAYER M4 ;
        RECT 536.104 105.032 536.256 105.184 ;
    END
    PORT
      LAYER M5 ;
        RECT 536.104 105.032 536.256 105.184 ;
    END
  END A1[10]

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
  END CE2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
  END CSB2

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.184 0.000 29.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.184 0.000 29.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.184 0.000 29.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.184 0.000 29.336 0.152 ;
    END
  END I2[0]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.488 0.000 29.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.488 0.000 29.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.488 0.000 29.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.488 0.000 29.640 0.152 ;
    END
  END I2[1]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.792 0.000 29.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.792 0.000 29.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.792 0.000 29.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.792 0.000 29.944 0.152 ;
    END
  END I2[2]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.096 0.000 30.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.096 0.000 30.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.096 0.000 30.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.096 0.000 30.248 0.152 ;
    END
  END I2[3]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
  END I2[4]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
  END I2[5]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
  END I2[6]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
  END I2[7]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
  END I2[8]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
  END I2[9]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
  END I2[10]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
  END I2[11]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
  END I2[12]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
  END I2[13]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
  END I2[14]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.984 0.000 52.136 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.984 0.000 52.136 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.984 0.000 52.136 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.984 0.000 52.136 0.152 ;
    END
  END I2[15]

  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
  END I2[16]

  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.672 0.000 58.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.672 0.000 58.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.672 0.000 58.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.672 0.000 58.824 0.152 ;
    END
  END I2[17]

  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
  END I2[18]

  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.280 0.000 59.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.280 0.000 59.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.280 0.000 59.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.280 0.000 59.432 0.152 ;
    END
  END I2[19]

  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
  END I2[20]

  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.968 0.000 66.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.968 0.000 66.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.968 0.000 66.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.968 0.000 66.120 0.152 ;
    END
  END I2[21]

  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.272 0.000 66.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.272 0.000 66.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.272 0.000 66.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.272 0.000 66.424 0.152 ;
    END
  END I2[22]

  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.576 0.000 66.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.576 0.000 66.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.576 0.000 66.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.576 0.000 66.728 0.152 ;
    END
  END I2[23]

  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.960 0.000 73.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.960 0.000 73.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.960 0.000 73.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.960 0.000 73.112 0.152 ;
    END
  END I2[24]

  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.264 0.000 73.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.264 0.000 73.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.264 0.000 73.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.264 0.000 73.416 0.152 ;
    END
  END I2[25]

  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.568 0.000 73.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.568 0.000 73.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.568 0.000 73.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.568 0.000 73.720 0.152 ;
    END
  END I2[26]

  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
  END I2[27]

  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
  END I2[28]

  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.560 0.000 80.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.560 0.000 80.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.560 0.000 80.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.560 0.000 80.712 0.152 ;
    END
  END I2[29]

  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.864 0.000 81.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.864 0.000 81.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.864 0.000 81.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.864 0.000 81.016 0.152 ;
    END
  END I2[30]

  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.168 0.000 81.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.168 0.000 81.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.168 0.000 81.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.168 0.000 81.320 0.152 ;
    END
  END I2[31]

  PIN I2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
  END I2[32]

  PIN I2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
  END I2[33]

  PIN I2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
  END I2[34]

  PIN I2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
  END I2[35]

  PIN I2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.848 0.000 95.000 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.848 0.000 95.000 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.848 0.000 95.000 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.848 0.000 95.000 0.152 ;
    END
  END I2[36]

  PIN I2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
  END I2[37]

  PIN I2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.456 0.000 95.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.456 0.000 95.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.456 0.000 95.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.456 0.000 95.608 0.152 ;
    END
  END I2[38]

  PIN I2[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.760 0.000 95.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.760 0.000 95.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.760 0.000 95.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.760 0.000 95.912 0.152 ;
    END
  END I2[39]

  PIN I2[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.144 0.000 102.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.144 0.000 102.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.144 0.000 102.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.144 0.000 102.296 0.152 ;
    END
  END I2[40]

  PIN I2[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.448 0.000 102.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.448 0.000 102.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.448 0.000 102.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.448 0.000 102.600 0.152 ;
    END
  END I2[41]

  PIN I2[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.752 0.000 102.904 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.752 0.000 102.904 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.752 0.000 102.904 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.752 0.000 102.904 0.152 ;
    END
  END I2[42]

  PIN I2[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.056 0.000 103.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.056 0.000 103.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.056 0.000 103.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.056 0.000 103.208 0.152 ;
    END
  END I2[43]

  PIN I2[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
  END I2[44]

  PIN I2[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
  END I2[45]

  PIN I2[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
  END I2[46]

  PIN I2[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
  END I2[47]

  PIN I2[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.736 0.000 116.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.736 0.000 116.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.736 0.000 116.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.736 0.000 116.888 0.152 ;
    END
  END I2[48]

  PIN I2[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.040 0.000 117.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 117.040 0.000 117.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 117.040 0.000 117.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.040 0.000 117.192 0.152 ;
    END
  END I2[49]

  PIN I2[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.344 0.000 117.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 117.344 0.000 117.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 117.344 0.000 117.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.344 0.000 117.496 0.152 ;
    END
  END I2[50]

  PIN I2[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.648 0.000 117.800 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 117.648 0.000 117.800 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 117.648 0.000 117.800 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.648 0.000 117.800 0.152 ;
    END
  END I2[51]

  PIN I2[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.032 0.000 124.184 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.032 0.000 124.184 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.032 0.000 124.184 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.032 0.000 124.184 0.152 ;
    END
  END I2[52]

  PIN I2[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.336 0.000 124.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.336 0.000 124.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.336 0.000 124.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.336 0.000 124.488 0.152 ;
    END
  END I2[53]

  PIN I2[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.640 0.000 124.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.640 0.000 124.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.640 0.000 124.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.640 0.000 124.792 0.152 ;
    END
  END I2[54]

  PIN I2[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.944 0.000 125.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.944 0.000 125.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.944 0.000 125.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.944 0.000 125.096 0.152 ;
    END
  END I2[55]

  PIN I2[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
  END I2[56]

  PIN I2[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.632 0.000 131.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.632 0.000 131.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.632 0.000 131.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.632 0.000 131.784 0.152 ;
    END
  END I2[57]

  PIN I2[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.936 0.000 132.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.936 0.000 132.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.936 0.000 132.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.936 0.000 132.088 0.152 ;
    END
  END I2[58]

  PIN I2[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.240 0.000 132.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.240 0.000 132.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.240 0.000 132.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 132.240 0.000 132.392 0.152 ;
    END
  END I2[59]

  PIN I2[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.624 0.000 138.776 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 138.624 0.000 138.776 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 138.624 0.000 138.776 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.624 0.000 138.776 0.152 ;
    END
  END I2[60]

  PIN I2[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.928 0.000 139.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 138.928 0.000 139.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 138.928 0.000 139.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.928 0.000 139.080 0.152 ;
    END
  END I2[61]

  PIN I2[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.232 0.000 139.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 139.232 0.000 139.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 139.232 0.000 139.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.232 0.000 139.384 0.152 ;
    END
  END I2[62]

  PIN I2[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.536 0.000 139.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 139.536 0.000 139.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 139.536 0.000 139.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.536 0.000 139.688 0.152 ;
    END
  END I2[63]

  PIN I2[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.920 0.000 146.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 145.920 0.000 146.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.920 0.000 146.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.920 0.000 146.072 0.152 ;
    END
  END I2[64]

  PIN I2[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
  END I2[65]

  PIN I2[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.528 0.000 146.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 146.528 0.000 146.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.528 0.000 146.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.528 0.000 146.680 0.152 ;
    END
  END I2[66]

  PIN I2[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.832 0.000 146.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 146.832 0.000 146.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.832 0.000 146.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.832 0.000 146.984 0.152 ;
    END
  END I2[67]

  PIN I2[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
  END I2[68]

  PIN I2[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
  END I2[69]

  PIN I2[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
  END I2[70]

  PIN I2[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
  END I2[71]

  PIN I2[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.512 0.000 160.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 160.512 0.000 160.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 160.512 0.000 160.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 160.512 0.000 160.664 0.152 ;
    END
  END I2[72]

  PIN I2[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.816 0.000 160.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 160.816 0.000 160.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 160.816 0.000 160.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 160.816 0.000 160.968 0.152 ;
    END
  END I2[73]

  PIN I2[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.120 0.000 161.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.120 0.000 161.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.120 0.000 161.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.120 0.000 161.272 0.152 ;
    END
  END I2[74]

  PIN I2[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.424 0.000 161.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.424 0.000 161.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.424 0.000 161.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.424 0.000 161.576 0.152 ;
    END
  END I2[75]

  PIN I2[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.808 0.000 167.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 167.808 0.000 167.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 167.808 0.000 167.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 167.808 0.000 167.960 0.152 ;
    END
  END I2[76]

  PIN I2[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.112 0.000 168.264 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 168.112 0.000 168.264 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 168.112 0.000 168.264 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 168.112 0.000 168.264 0.152 ;
    END
  END I2[77]

  PIN I2[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.416 0.000 168.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 168.416 0.000 168.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 168.416 0.000 168.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 168.416 0.000 168.568 0.152 ;
    END
  END I2[78]

  PIN I2[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.720 0.000 168.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 168.720 0.000 168.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 168.720 0.000 168.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 168.720 0.000 168.872 0.152 ;
    END
  END I2[79]

  PIN I2[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
  END I2[80]

  PIN I2[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
  END I2[81]

  PIN I2[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
  END I2[82]

  PIN I2[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
  END I2[83]

  PIN I2[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.400 0.000 182.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 182.400 0.000 182.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 182.400 0.000 182.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 182.400 0.000 182.552 0.152 ;
    END
  END I2[84]

  PIN I2[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.704 0.000 182.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 182.704 0.000 182.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 182.704 0.000 182.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 182.704 0.000 182.856 0.152 ;
    END
  END I2[85]

  PIN I2[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.008 0.000 183.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 183.008 0.000 183.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 183.008 0.000 183.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 183.008 0.000 183.160 0.152 ;
    END
  END I2[86]

  PIN I2[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.312 0.000 183.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 183.312 0.000 183.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 183.312 0.000 183.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 183.312 0.000 183.464 0.152 ;
    END
  END I2[87]

  PIN I2[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.696 0.000 189.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 189.696 0.000 189.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 189.696 0.000 189.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 189.696 0.000 189.848 0.152 ;
    END
  END I2[88]

  PIN I2[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.000 0.000 190.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.000 0.000 190.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.000 0.000 190.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.000 0.000 190.152 0.152 ;
    END
  END I2[89]

  PIN I2[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.304 0.000 190.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.304 0.000 190.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.304 0.000 190.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.304 0.000 190.456 0.152 ;
    END
  END I2[90]

  PIN I2[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
  END I2[91]

  PIN I2[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.992 0.000 197.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 196.992 0.000 197.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 196.992 0.000 197.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 196.992 0.000 197.144 0.152 ;
    END
  END I2[92]

  PIN I2[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.296 0.000 197.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.296 0.000 197.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.296 0.000 197.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 197.296 0.000 197.448 0.152 ;
    END
  END I2[93]

  PIN I2[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.600 0.000 197.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.600 0.000 197.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.600 0.000 197.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 197.600 0.000 197.752 0.152 ;
    END
  END I2[94]

  PIN I2[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.904 0.000 198.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.904 0.000 198.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.904 0.000 198.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 197.904 0.000 198.056 0.152 ;
    END
  END I2[95]

  PIN I2[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.288 0.000 204.440 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 204.288 0.000 204.440 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 204.288 0.000 204.440 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 204.288 0.000 204.440 0.152 ;
    END
  END I2[96]

  PIN I2[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.592 0.000 204.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 204.592 0.000 204.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 204.592 0.000 204.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 204.592 0.000 204.744 0.152 ;
    END
  END I2[97]

  PIN I2[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.896 0.000 205.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 204.896 0.000 205.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 204.896 0.000 205.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 204.896 0.000 205.048 0.152 ;
    END
  END I2[98]

  PIN I2[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.200 0.000 205.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.200 0.000 205.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.200 0.000 205.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.200 0.000 205.352 0.152 ;
    END
  END I2[99]

  PIN I2[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.584 0.000 211.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 211.584 0.000 211.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 211.584 0.000 211.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 211.584 0.000 211.736 0.152 ;
    END
  END I2[100]

  PIN I2[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.888 0.000 212.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 211.888 0.000 212.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 211.888 0.000 212.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 211.888 0.000 212.040 0.152 ;
    END
  END I2[101]

  PIN I2[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.192 0.000 212.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 212.192 0.000 212.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 212.192 0.000 212.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 212.192 0.000 212.344 0.152 ;
    END
  END I2[102]

  PIN I2[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.496 0.000 212.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 212.496 0.000 212.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 212.496 0.000 212.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 212.496 0.000 212.648 0.152 ;
    END
  END I2[103]

  PIN I2[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.880 0.000 219.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 218.880 0.000 219.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 218.880 0.000 219.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 218.880 0.000 219.032 0.152 ;
    END
  END I2[104]

  PIN I2[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.184 0.000 219.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 219.184 0.000 219.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 219.184 0.000 219.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 219.184 0.000 219.336 0.152 ;
    END
  END I2[105]

  PIN I2[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.488 0.000 219.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 219.488 0.000 219.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 219.488 0.000 219.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 219.488 0.000 219.640 0.152 ;
    END
  END I2[106]

  PIN I2[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.792 0.000 219.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 219.792 0.000 219.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 219.792 0.000 219.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 219.792 0.000 219.944 0.152 ;
    END
  END I2[107]

  PIN I2[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.176 0.000 226.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 226.176 0.000 226.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 226.176 0.000 226.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 226.176 0.000 226.328 0.152 ;
    END
  END I2[108]

  PIN I2[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.480 0.000 226.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 226.480 0.000 226.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 226.480 0.000 226.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 226.480 0.000 226.632 0.152 ;
    END
  END I2[109]

  PIN I2[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.784 0.000 226.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 226.784 0.000 226.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 226.784 0.000 226.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 226.784 0.000 226.936 0.152 ;
    END
  END I2[110]

  PIN I2[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 227.088 0.000 227.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 227.088 0.000 227.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 227.088 0.000 227.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 227.088 0.000 227.240 0.152 ;
    END
  END I2[111]

  PIN I2[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 233.472 0.000 233.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 233.472 0.000 233.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 233.472 0.000 233.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 233.472 0.000 233.624 0.152 ;
    END
  END I2[112]

  PIN I2[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 233.776 0.000 233.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 233.776 0.000 233.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 233.776 0.000 233.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 233.776 0.000 233.928 0.152 ;
    END
  END I2[113]

  PIN I2[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.080 0.000 234.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 234.080 0.000 234.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 234.080 0.000 234.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 234.080 0.000 234.232 0.152 ;
    END
  END I2[114]

  PIN I2[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.384 0.000 234.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 234.384 0.000 234.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 234.384 0.000 234.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 234.384 0.000 234.536 0.152 ;
    END
  END I2[115]

  PIN I2[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 240.768 0.000 240.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 240.768 0.000 240.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 240.768 0.000 240.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 240.768 0.000 240.920 0.152 ;
    END
  END I2[116]

  PIN I2[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.072 0.000 241.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 241.072 0.000 241.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 241.072 0.000 241.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 241.072 0.000 241.224 0.152 ;
    END
  END I2[117]

  PIN I2[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.376 0.000 241.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 241.376 0.000 241.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 241.376 0.000 241.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 241.376 0.000 241.528 0.152 ;
    END
  END I2[118]

  PIN I2[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.680 0.000 241.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 241.680 0.000 241.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 241.680 0.000 241.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 241.680 0.000 241.832 0.152 ;
    END
  END I2[119]

  PIN I2[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.064 0.000 248.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 248.064 0.000 248.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 248.064 0.000 248.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 248.064 0.000 248.216 0.152 ;
    END
  END I2[120]

  PIN I2[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.368 0.000 248.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 248.368 0.000 248.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 248.368 0.000 248.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 248.368 0.000 248.520 0.152 ;
    END
  END I2[121]

  PIN I2[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.672 0.000 248.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 248.672 0.000 248.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 248.672 0.000 248.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 248.672 0.000 248.824 0.152 ;
    END
  END I2[122]

  PIN I2[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.976 0.000 249.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 248.976 0.000 249.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 248.976 0.000 249.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 248.976 0.000 249.128 0.152 ;
    END
  END I2[123]

  PIN I2[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.360 0.000 255.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 255.360 0.000 255.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 255.360 0.000 255.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 255.360 0.000 255.512 0.152 ;
    END
  END I2[124]

  PIN I2[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.664 0.000 255.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 255.664 0.000 255.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 255.664 0.000 255.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 255.664 0.000 255.816 0.152 ;
    END
  END I2[125]

  PIN I2[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.968 0.000 256.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 255.968 0.000 256.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 255.968 0.000 256.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 255.968 0.000 256.120 0.152 ;
    END
  END I2[126]

  PIN I2[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 256.272 0.000 256.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 256.272 0.000 256.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 256.272 0.000 256.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 256.272 0.000 256.424 0.152 ;
    END
  END I2[127]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 141.512 0.152 141.664 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 141.512 0.152 141.664 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 141.512 0.152 141.664 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 141.512 0.152 141.664 ;
    END
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 137.864 0.152 138.016 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 137.864 0.152 138.016 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 137.864 0.152 138.016 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 137.864 0.152 138.016 ;
    END
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 134.216 0.152 134.368 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 134.216 0.152 134.368 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 134.216 0.152 134.368 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 134.216 0.152 134.368 ;
    END
  END A2[2]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 130.568 0.152 130.720 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 130.568 0.152 130.720 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 130.568 0.152 130.720 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 130.568 0.152 130.720 ;
    END
  END A2[3]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 126.920 0.152 127.072 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 126.920 0.152 127.072 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 126.920 0.152 127.072 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 126.920 0.152 127.072 ;
    END
  END A2[4]

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 123.272 0.152 123.424 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 123.272 0.152 123.424 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 123.272 0.152 123.424 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 123.272 0.152 123.424 ;
    END
  END A2[5]

  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 119.624 0.152 119.776 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 119.624 0.152 119.776 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 119.624 0.152 119.776 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 119.624 0.152 119.776 ;
    END
  END A2[6]

  PIN A2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 115.976 0.152 116.128 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 115.976 0.152 116.128 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 115.976 0.152 116.128 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 115.976 0.152 116.128 ;
    END
  END A2[7]

  PIN A2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 112.328 0.152 112.480 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 112.328 0.152 112.480 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 112.328 0.152 112.480 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 112.328 0.152 112.480 ;
    END
  END A2[8]

  PIN A2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 108.680 0.152 108.832 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 108.680 0.152 108.832 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 108.680 0.152 108.832 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 108.680 0.152 108.832 ;
    END
  END A2[9]

  PIN A2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 105.032 0.152 105.184 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 105.032 0.152 105.184 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 105.032 0.152 105.184 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 105.032 0.152 105.184 ;
    END
  END A2[10]

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 40.432 0.152 40.584 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 40.432 0.152 40.584 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 40.432 0.152 40.584 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 40.432 0.152 40.584 ;
    END
  END WEB2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 5.195 159.728 7.195 161.728 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.195 159.728 7.195 161.728 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.195 159.728 7.195 161.728 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 7.915 159.728 9.915 161.728 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.915 159.728 9.915 161.728 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.915 159.728 9.915 161.728 ;
    END
  END VSS

  OBS
    LAYER M2 ;
      RECT 520.144 0.000 536.256 0.304 ;
      RECT 513.760 0.000 519.688 0.304 ;
      RECT 507.376 0.000 513.304 0.304 ;
      RECT 500.992 0.000 506.920 0.304 ;
      RECT 493.696 0.000 499.624 0.304 ;
      RECT 486.400 0.000 492.328 0.304 ;
      RECT 479.104 0.000 485.032 0.304 ;
      RECT 471.808 0.000 477.736 0.304 ;
      RECT 464.512 0.000 470.440 0.304 ;
      RECT 457.216 0.000 463.144 0.304 ;
      RECT 449.920 0.000 455.848 0.304 ;
      RECT 442.624 0.000 448.552 0.304 ;
      RECT 435.328 0.000 441.256 0.304 ;
      RECT 428.032 0.000 433.960 0.304 ;
      RECT 420.736 0.000 426.664 0.304 ;
      RECT 413.440 0.000 419.368 0.304 ;
      RECT 406.144 0.000 412.072 0.304 ;
      RECT 398.848 0.000 404.776 0.304 ;
      RECT 391.552 0.000 397.480 0.304 ;
      RECT 384.256 0.000 390.184 0.304 ;
      RECT 376.960 0.000 382.888 0.304 ;
      RECT 369.664 0.000 375.592 0.304 ;
      RECT 362.368 0.000 368.296 0.304 ;
      RECT 355.072 0.000 361.000 0.304 ;
      RECT 347.776 0.000 353.704 0.304 ;
      RECT 340.480 0.000 346.408 0.304 ;
      RECT 333.184 0.000 339.112 0.304 ;
      RECT 325.888 0.000 331.816 0.304 ;
      RECT 318.592 0.000 324.520 0.304 ;
      RECT 311.296 0.000 317.224 0.304 ;
      RECT 304.000 0.000 309.928 0.304 ;
      RECT 296.704 0.000 302.632 0.304 ;
      RECT 289.408 0.000 295.336 0.304 ;
      RECT 282.112 0.000 288.040 0.304 ;
      RECT 274.816 0.000 280.744 0.304 ;
      RECT 535.952 141.816 536.256 159.576 ;
      RECT 535.952 138.168 536.256 141.360 ;
      RECT 535.952 134.520 536.256 137.712 ;
      RECT 535.952 130.872 536.256 134.064 ;
      RECT 535.952 127.224 536.256 130.416 ;
      RECT 535.952 123.576 536.256 126.768 ;
      RECT 535.952 119.928 536.256 123.120 ;
      RECT 535.952 116.280 536.256 119.472 ;
      RECT 535.952 112.632 536.256 115.824 ;
      RECT 535.952 108.984 536.256 112.176 ;
      RECT 535.952 105.336 536.256 108.528 ;
      RECT 535.952 40.736 536.256 104.880 ;
      RECT 535.952 0.304 536.256 40.280 ;
      RECT 0.000 0.000 16.264 0.304 ;
      RECT 16.720 0.000 22.648 0.304 ;
      RECT 23.104 0.000 29.032 0.304 ;
      RECT 30.400 0.000 36.328 0.304 ;
      RECT 37.696 0.000 43.624 0.304 ;
      RECT 44.992 0.000 50.920 0.304 ;
      RECT 52.288 0.000 58.216 0.304 ;
      RECT 59.584 0.000 65.512 0.304 ;
      RECT 66.880 0.000 72.808 0.304 ;
      RECT 74.176 0.000 80.104 0.304 ;
      RECT 81.472 0.000 87.400 0.304 ;
      RECT 88.768 0.000 94.696 0.304 ;
      RECT 96.064 0.000 101.992 0.304 ;
      RECT 103.360 0.000 109.288 0.304 ;
      RECT 110.656 0.000 116.584 0.304 ;
      RECT 117.952 0.000 123.880 0.304 ;
      RECT 125.248 0.000 131.176 0.304 ;
      RECT 132.544 0.000 138.472 0.304 ;
      RECT 139.840 0.000 145.768 0.304 ;
      RECT 147.136 0.000 153.064 0.304 ;
      RECT 154.432 0.000 160.360 0.304 ;
      RECT 161.728 0.000 167.656 0.304 ;
      RECT 169.024 0.000 174.952 0.304 ;
      RECT 176.320 0.000 182.248 0.304 ;
      RECT 183.616 0.000 189.544 0.304 ;
      RECT 190.912 0.000 196.840 0.304 ;
      RECT 198.208 0.000 204.136 0.304 ;
      RECT 205.504 0.000 211.432 0.304 ;
      RECT 212.800 0.000 218.728 0.304 ;
      RECT 220.096 0.000 226.024 0.304 ;
      RECT 227.392 0.000 233.320 0.304 ;
      RECT 234.688 0.000 240.616 0.304 ;
      RECT 241.984 0.000 247.912 0.304 ;
      RECT 249.280 0.000 255.208 0.304 ;
      RECT 256.576 0.000 273.448 0.304 ;
      RECT 0.000 141.816 0.304 159.576 ;
      RECT 0.000 138.168 0.304 141.360 ;
      RECT 0.000 134.520 0.304 137.712 ;
      RECT 0.000 130.872 0.304 134.064 ;
      RECT 0.000 127.224 0.304 130.416 ;
      RECT 0.000 123.576 0.304 126.768 ;
      RECT 0.000 119.928 0.304 123.120 ;
      RECT 0.000 116.280 0.304 119.472 ;
      RECT 0.000 112.632 0.304 115.824 ;
      RECT 0.000 108.984 0.304 112.176 ;
      RECT 0.000 105.336 0.304 108.528 ;
      RECT 0.000 40.736 0.304 104.880 ;
      RECT 0.000 0.304 0.304 40.280 ;
      RECT 0.000 159.576 5.043 161.728 ;
      RECT 7.355 159.576 7.763 161.728 ;
      RECT 10.067 159.576 536.256 161.728 ;
      RECT 0.304 0.304 535.952 159.576 ;
    LAYER M3 ;
      RECT 520.144 0.000 536.256 0.304 ;
      RECT 513.760 0.000 519.688 0.304 ;
      RECT 507.376 0.000 513.304 0.304 ;
      RECT 500.992 0.000 506.920 0.304 ;
      RECT 493.696 0.000 499.624 0.304 ;
      RECT 486.400 0.000 492.328 0.304 ;
      RECT 479.104 0.000 485.032 0.304 ;
      RECT 471.808 0.000 477.736 0.304 ;
      RECT 464.512 0.000 470.440 0.304 ;
      RECT 457.216 0.000 463.144 0.304 ;
      RECT 449.920 0.000 455.848 0.304 ;
      RECT 442.624 0.000 448.552 0.304 ;
      RECT 435.328 0.000 441.256 0.304 ;
      RECT 428.032 0.000 433.960 0.304 ;
      RECT 420.736 0.000 426.664 0.304 ;
      RECT 413.440 0.000 419.368 0.304 ;
      RECT 406.144 0.000 412.072 0.304 ;
      RECT 398.848 0.000 404.776 0.304 ;
      RECT 391.552 0.000 397.480 0.304 ;
      RECT 384.256 0.000 390.184 0.304 ;
      RECT 376.960 0.000 382.888 0.304 ;
      RECT 369.664 0.000 375.592 0.304 ;
      RECT 362.368 0.000 368.296 0.304 ;
      RECT 355.072 0.000 361.000 0.304 ;
      RECT 347.776 0.000 353.704 0.304 ;
      RECT 340.480 0.000 346.408 0.304 ;
      RECT 333.184 0.000 339.112 0.304 ;
      RECT 325.888 0.000 331.816 0.304 ;
      RECT 318.592 0.000 324.520 0.304 ;
      RECT 311.296 0.000 317.224 0.304 ;
      RECT 304.000 0.000 309.928 0.304 ;
      RECT 296.704 0.000 302.632 0.304 ;
      RECT 289.408 0.000 295.336 0.304 ;
      RECT 282.112 0.000 288.040 0.304 ;
      RECT 274.816 0.000 280.744 0.304 ;
      RECT 535.952 141.816 536.256 159.576 ;
      RECT 535.952 138.168 536.256 141.360 ;
      RECT 535.952 134.520 536.256 137.712 ;
      RECT 535.952 130.872 536.256 134.064 ;
      RECT 535.952 127.224 536.256 130.416 ;
      RECT 535.952 123.576 536.256 126.768 ;
      RECT 535.952 119.928 536.256 123.120 ;
      RECT 535.952 116.280 536.256 119.472 ;
      RECT 535.952 112.632 536.256 115.824 ;
      RECT 535.952 108.984 536.256 112.176 ;
      RECT 535.952 105.336 536.256 108.528 ;
      RECT 535.952 40.736 536.256 104.880 ;
      RECT 535.952 0.304 536.256 40.280 ;
      RECT 0.000 0.000 16.264 0.304 ;
      RECT 16.720 0.000 22.648 0.304 ;
      RECT 23.104 0.000 29.032 0.304 ;
      RECT 30.400 0.000 36.328 0.304 ;
      RECT 37.696 0.000 43.624 0.304 ;
      RECT 44.992 0.000 50.920 0.304 ;
      RECT 52.288 0.000 58.216 0.304 ;
      RECT 59.584 0.000 65.512 0.304 ;
      RECT 66.880 0.000 72.808 0.304 ;
      RECT 74.176 0.000 80.104 0.304 ;
      RECT 81.472 0.000 87.400 0.304 ;
      RECT 88.768 0.000 94.696 0.304 ;
      RECT 96.064 0.000 101.992 0.304 ;
      RECT 103.360 0.000 109.288 0.304 ;
      RECT 110.656 0.000 116.584 0.304 ;
      RECT 117.952 0.000 123.880 0.304 ;
      RECT 125.248 0.000 131.176 0.304 ;
      RECT 132.544 0.000 138.472 0.304 ;
      RECT 139.840 0.000 145.768 0.304 ;
      RECT 147.136 0.000 153.064 0.304 ;
      RECT 154.432 0.000 160.360 0.304 ;
      RECT 161.728 0.000 167.656 0.304 ;
      RECT 169.024 0.000 174.952 0.304 ;
      RECT 176.320 0.000 182.248 0.304 ;
      RECT 183.616 0.000 189.544 0.304 ;
      RECT 190.912 0.000 196.840 0.304 ;
      RECT 198.208 0.000 204.136 0.304 ;
      RECT 205.504 0.000 211.432 0.304 ;
      RECT 212.800 0.000 218.728 0.304 ;
      RECT 220.096 0.000 226.024 0.304 ;
      RECT 227.392 0.000 233.320 0.304 ;
      RECT 234.688 0.000 240.616 0.304 ;
      RECT 241.984 0.000 247.912 0.304 ;
      RECT 249.280 0.000 255.208 0.304 ;
      RECT 256.576 0.000 273.448 0.304 ;
      RECT 0.000 141.816 0.304 159.576 ;
      RECT 0.000 138.168 0.304 141.360 ;
      RECT 0.000 134.520 0.304 137.712 ;
      RECT 0.000 130.872 0.304 134.064 ;
      RECT 0.000 127.224 0.304 130.416 ;
      RECT 0.000 123.576 0.304 126.768 ;
      RECT 0.000 119.928 0.304 123.120 ;
      RECT 0.000 116.280 0.304 119.472 ;
      RECT 0.000 112.632 0.304 115.824 ;
      RECT 0.000 108.984 0.304 112.176 ;
      RECT 0.000 105.336 0.304 108.528 ;
      RECT 0.000 40.736 0.304 104.880 ;
      RECT 0.000 0.304 0.304 40.280 ;
      RECT 0.000 159.576 5.043 161.728 ;
      RECT 7.355 159.576 7.763 161.728 ;
      RECT 10.067 159.576 536.256 161.728 ;
      RECT 0.304 0.304 535.952 159.576 ;
    LAYER M4 ;
      RECT 520.144 0.000 536.256 0.304 ;
      RECT 513.760 0.000 519.688 0.304 ;
      RECT 507.376 0.000 513.304 0.304 ;
      RECT 500.992 0.000 506.920 0.304 ;
      RECT 493.696 0.000 499.624 0.304 ;
      RECT 486.400 0.000 492.328 0.304 ;
      RECT 479.104 0.000 485.032 0.304 ;
      RECT 471.808 0.000 477.736 0.304 ;
      RECT 464.512 0.000 470.440 0.304 ;
      RECT 457.216 0.000 463.144 0.304 ;
      RECT 449.920 0.000 455.848 0.304 ;
      RECT 442.624 0.000 448.552 0.304 ;
      RECT 435.328 0.000 441.256 0.304 ;
      RECT 428.032 0.000 433.960 0.304 ;
      RECT 420.736 0.000 426.664 0.304 ;
      RECT 413.440 0.000 419.368 0.304 ;
      RECT 406.144 0.000 412.072 0.304 ;
      RECT 398.848 0.000 404.776 0.304 ;
      RECT 391.552 0.000 397.480 0.304 ;
      RECT 384.256 0.000 390.184 0.304 ;
      RECT 376.960 0.000 382.888 0.304 ;
      RECT 369.664 0.000 375.592 0.304 ;
      RECT 362.368 0.000 368.296 0.304 ;
      RECT 355.072 0.000 361.000 0.304 ;
      RECT 347.776 0.000 353.704 0.304 ;
      RECT 340.480 0.000 346.408 0.304 ;
      RECT 333.184 0.000 339.112 0.304 ;
      RECT 325.888 0.000 331.816 0.304 ;
      RECT 318.592 0.000 324.520 0.304 ;
      RECT 311.296 0.000 317.224 0.304 ;
      RECT 304.000 0.000 309.928 0.304 ;
      RECT 296.704 0.000 302.632 0.304 ;
      RECT 289.408 0.000 295.336 0.304 ;
      RECT 282.112 0.000 288.040 0.304 ;
      RECT 274.816 0.000 280.744 0.304 ;
      RECT 535.952 141.816 536.256 159.576 ;
      RECT 535.952 138.168 536.256 141.360 ;
      RECT 535.952 134.520 536.256 137.712 ;
      RECT 535.952 130.872 536.256 134.064 ;
      RECT 535.952 127.224 536.256 130.416 ;
      RECT 535.952 123.576 536.256 126.768 ;
      RECT 535.952 119.928 536.256 123.120 ;
      RECT 535.952 116.280 536.256 119.472 ;
      RECT 535.952 112.632 536.256 115.824 ;
      RECT 535.952 108.984 536.256 112.176 ;
      RECT 535.952 105.336 536.256 108.528 ;
      RECT 535.952 40.736 536.256 104.880 ;
      RECT 535.952 0.304 536.256 40.280 ;
      RECT 0.000 0.000 16.264 0.304 ;
      RECT 16.720 0.000 22.648 0.304 ;
      RECT 23.104 0.000 29.032 0.304 ;
      RECT 30.400 0.000 36.328 0.304 ;
      RECT 37.696 0.000 43.624 0.304 ;
      RECT 44.992 0.000 50.920 0.304 ;
      RECT 52.288 0.000 58.216 0.304 ;
      RECT 59.584 0.000 65.512 0.304 ;
      RECT 66.880 0.000 72.808 0.304 ;
      RECT 74.176 0.000 80.104 0.304 ;
      RECT 81.472 0.000 87.400 0.304 ;
      RECT 88.768 0.000 94.696 0.304 ;
      RECT 96.064 0.000 101.992 0.304 ;
      RECT 103.360 0.000 109.288 0.304 ;
      RECT 110.656 0.000 116.584 0.304 ;
      RECT 117.952 0.000 123.880 0.304 ;
      RECT 125.248 0.000 131.176 0.304 ;
      RECT 132.544 0.000 138.472 0.304 ;
      RECT 139.840 0.000 145.768 0.304 ;
      RECT 147.136 0.000 153.064 0.304 ;
      RECT 154.432 0.000 160.360 0.304 ;
      RECT 161.728 0.000 167.656 0.304 ;
      RECT 169.024 0.000 174.952 0.304 ;
      RECT 176.320 0.000 182.248 0.304 ;
      RECT 183.616 0.000 189.544 0.304 ;
      RECT 190.912 0.000 196.840 0.304 ;
      RECT 198.208 0.000 204.136 0.304 ;
      RECT 205.504 0.000 211.432 0.304 ;
      RECT 212.800 0.000 218.728 0.304 ;
      RECT 220.096 0.000 226.024 0.304 ;
      RECT 227.392 0.000 233.320 0.304 ;
      RECT 234.688 0.000 240.616 0.304 ;
      RECT 241.984 0.000 247.912 0.304 ;
      RECT 249.280 0.000 255.208 0.304 ;
      RECT 256.576 0.000 273.448 0.304 ;
      RECT 0.000 141.816 0.304 159.576 ;
      RECT 0.000 138.168 0.304 141.360 ;
      RECT 0.000 134.520 0.304 137.712 ;
      RECT 0.000 130.872 0.304 134.064 ;
      RECT 0.000 127.224 0.304 130.416 ;
      RECT 0.000 123.576 0.304 126.768 ;
      RECT 0.000 119.928 0.304 123.120 ;
      RECT 0.000 116.280 0.304 119.472 ;
      RECT 0.000 112.632 0.304 115.824 ;
      RECT 0.000 108.984 0.304 112.176 ;
      RECT 0.000 105.336 0.304 108.528 ;
      RECT 0.000 40.736 0.304 104.880 ;
      RECT 0.000 0.304 0.304 40.280 ;
      RECT 0.000 159.576 5.043 161.728 ;
      RECT 7.355 159.576 7.763 161.728 ;
      RECT 10.067 159.576 536.256 161.728 ;
      RECT 0.304 0.304 535.952 159.576 ;
    LAYER M5 ;
      RECT 520.144 0.000 536.256 0.304 ;
      RECT 513.760 0.000 519.688 0.304 ;
      RECT 507.376 0.000 513.304 0.304 ;
      RECT 500.992 0.000 506.920 0.304 ;
      RECT 493.696 0.000 499.624 0.304 ;
      RECT 486.400 0.000 492.328 0.304 ;
      RECT 479.104 0.000 485.032 0.304 ;
      RECT 471.808 0.000 477.736 0.304 ;
      RECT 464.512 0.000 470.440 0.304 ;
      RECT 457.216 0.000 463.144 0.304 ;
      RECT 449.920 0.000 455.848 0.304 ;
      RECT 442.624 0.000 448.552 0.304 ;
      RECT 435.328 0.000 441.256 0.304 ;
      RECT 428.032 0.000 433.960 0.304 ;
      RECT 420.736 0.000 426.664 0.304 ;
      RECT 413.440 0.000 419.368 0.304 ;
      RECT 406.144 0.000 412.072 0.304 ;
      RECT 398.848 0.000 404.776 0.304 ;
      RECT 391.552 0.000 397.480 0.304 ;
      RECT 384.256 0.000 390.184 0.304 ;
      RECT 376.960 0.000 382.888 0.304 ;
      RECT 369.664 0.000 375.592 0.304 ;
      RECT 362.368 0.000 368.296 0.304 ;
      RECT 355.072 0.000 361.000 0.304 ;
      RECT 347.776 0.000 353.704 0.304 ;
      RECT 340.480 0.000 346.408 0.304 ;
      RECT 333.184 0.000 339.112 0.304 ;
      RECT 325.888 0.000 331.816 0.304 ;
      RECT 318.592 0.000 324.520 0.304 ;
      RECT 311.296 0.000 317.224 0.304 ;
      RECT 304.000 0.000 309.928 0.304 ;
      RECT 296.704 0.000 302.632 0.304 ;
      RECT 289.408 0.000 295.336 0.304 ;
      RECT 282.112 0.000 288.040 0.304 ;
      RECT 274.816 0.000 280.744 0.304 ;
      RECT 535.952 141.816 536.256 159.576 ;
      RECT 535.952 138.168 536.256 141.360 ;
      RECT 535.952 134.520 536.256 137.712 ;
      RECT 535.952 130.872 536.256 134.064 ;
      RECT 535.952 127.224 536.256 130.416 ;
      RECT 535.952 123.576 536.256 126.768 ;
      RECT 535.952 119.928 536.256 123.120 ;
      RECT 535.952 116.280 536.256 119.472 ;
      RECT 535.952 112.632 536.256 115.824 ;
      RECT 535.952 108.984 536.256 112.176 ;
      RECT 535.952 105.336 536.256 108.528 ;
      RECT 535.952 40.736 536.256 104.880 ;
      RECT 535.952 0.304 536.256 40.280 ;
      RECT 0.000 0.000 16.264 0.304 ;
      RECT 16.720 0.000 22.648 0.304 ;
      RECT 23.104 0.000 29.032 0.304 ;
      RECT 30.400 0.000 36.328 0.304 ;
      RECT 37.696 0.000 43.624 0.304 ;
      RECT 44.992 0.000 50.920 0.304 ;
      RECT 52.288 0.000 58.216 0.304 ;
      RECT 59.584 0.000 65.512 0.304 ;
      RECT 66.880 0.000 72.808 0.304 ;
      RECT 74.176 0.000 80.104 0.304 ;
      RECT 81.472 0.000 87.400 0.304 ;
      RECT 88.768 0.000 94.696 0.304 ;
      RECT 96.064 0.000 101.992 0.304 ;
      RECT 103.360 0.000 109.288 0.304 ;
      RECT 110.656 0.000 116.584 0.304 ;
      RECT 117.952 0.000 123.880 0.304 ;
      RECT 125.248 0.000 131.176 0.304 ;
      RECT 132.544 0.000 138.472 0.304 ;
      RECT 139.840 0.000 145.768 0.304 ;
      RECT 147.136 0.000 153.064 0.304 ;
      RECT 154.432 0.000 160.360 0.304 ;
      RECT 161.728 0.000 167.656 0.304 ;
      RECT 169.024 0.000 174.952 0.304 ;
      RECT 176.320 0.000 182.248 0.304 ;
      RECT 183.616 0.000 189.544 0.304 ;
      RECT 190.912 0.000 196.840 0.304 ;
      RECT 198.208 0.000 204.136 0.304 ;
      RECT 205.504 0.000 211.432 0.304 ;
      RECT 212.800 0.000 218.728 0.304 ;
      RECT 220.096 0.000 226.024 0.304 ;
      RECT 227.392 0.000 233.320 0.304 ;
      RECT 234.688 0.000 240.616 0.304 ;
      RECT 241.984 0.000 247.912 0.304 ;
      RECT 249.280 0.000 255.208 0.304 ;
      RECT 256.576 0.000 273.448 0.304 ;
      RECT 0.000 141.816 0.304 159.576 ;
      RECT 0.000 138.168 0.304 141.360 ;
      RECT 0.000 134.520 0.304 137.712 ;
      RECT 0.000 130.872 0.304 134.064 ;
      RECT 0.000 127.224 0.304 130.416 ;
      RECT 0.000 123.576 0.304 126.768 ;
      RECT 0.000 119.928 0.304 123.120 ;
      RECT 0.000 116.280 0.304 119.472 ;
      RECT 0.000 112.632 0.304 115.824 ;
      RECT 0.000 108.984 0.304 112.176 ;
      RECT 0.000 105.336 0.304 108.528 ;
      RECT 0.000 40.736 0.304 104.880 ;
      RECT 0.000 0.304 0.304 40.280 ;
      RECT 0.000 159.576 5.043 161.728 ;
      RECT 7.355 159.576 7.763 161.728 ;
      RECT 10.067 159.576 536.256 161.728 ;
      RECT 0.304 0.304 535.952 159.576 ;
  END

END SRAM_128x1296_2P

END LIBRARY
