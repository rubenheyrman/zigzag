
//------> /esat/micas-data/software/Mentor/catapult_10.5c/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /esat/micas-data/software/Mentor/catapult_10.5c/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> ../td_ccore_solutions/O_addr_cnt_5_O_addr_type_L1_1__7448a59bcc55848f49259c21df88d8bc12ff1_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   r0678912@amazone.esat.kuleuven.be
//  Generated date: Tue Jul 13 10:58:06 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    O_addr_cnt_5_O_addr_type_L1_1
// ------------------------------------------------------------------


module O_addr_cnt_5_O_addr_type_L1_1 (
  loop_bound, tile_sizes, pntr_in, pntr_out, irrel_at_max_out, irrel_at_zero_out,
      all_at_max_1_out, counter_in, counter_out, tile_bound_in, tile_bound_out
);
  input [24:0] loop_bound;
  input [24:0] tile_sizes;
  input [4:0] pntr_in;
  output [4:0] pntr_out;
  output irrel_at_max_out;
  output irrel_at_zero_out;
  output all_at_max_1_out;
  input [24:0] counter_in;
  output [24:0] counter_out;
  input [24:0] tile_bound_in;
  output [24:0] tile_bound_out;


  // Interconnect Declarations
  wire for_1_unequal_4_tmp;
  wire [5:0] operator_5_false_acc_4_tmp;
  wire [6:0] nl_operator_5_false_acc_4_tmp;
  wire for_1_unequal_3_tmp;
  wire [5:0] operator_5_false_acc_3_tmp;
  wire [6:0] nl_operator_5_false_acc_3_tmp;
  wire for_1_unequal_2_tmp;
  wire [5:0] operator_5_false_acc_2_tmp;
  wire [6:0] nl_operator_5_false_acc_2_tmp;
  wire for_1_unequal_1_tmp;
  wire [5:0] operator_5_false_acc_1_tmp;
  wire [6:0] nl_operator_5_false_acc_1_tmp;
  wire for_1_for_1_for_1_for_1_nor_tmp;
  wire and_dcpl;
  wire and_dcpl_3;
  wire and_dcpl_4;
  wire and_dcpl_9;
  wire and_dcpl_10;
  wire and_dcpl_12;
  wire or_tmp_4;
  wire and_tmp;
  wire and_dcpl_24;
  wire or_tmp_14;
  wire mux_tmp_24;
  wire mux_tmp_25;
  wire and_dcpl_27;
  wire and_dcpl_28;
  wire or_dcpl_10;
  wire or_tmp_31;
  wire mux_tmp_30;
  wire and_dcpl_35;
  wire or_dcpl_13;
  wire or_tmp_41;
  wire not_tmp_24;
  wire and_dcpl_38;
  wire and_dcpl_46;
  wire or_dcpl_16;
  wire or_dcpl_18;
  wire or_dcpl_21;
  wire and_dcpl_53;
  wire or_dcpl_23;
  wire or_dcpl_25;
  wire or_tmp_48;
  wire and_dcpl_64;
  wire and_dcpl_65;
  wire [4:0] counter_buf_4_1_mx0;
  wire [4:0] counter_buf_3_1_mx0;
  wire [4:0] counter_buf_2_1_mx0;
  wire [4:0] counter_buf_1_1_mx0;
  wire equal_mdf_1;
  wire [5:0] operator_5_false_acc_cse_1;
  wire [6:0] nl_operator_5_false_acc_cse_1;
  wire [4:0] counter_buf_0_1_mx1;
  wire mux_9_cse;
  wire or_89_cse;
  wire or_79_cse;
  wire or_75_cse;
  wire or_82_cse;
  wire or_20_cse;
  wire nor_16_cse;
  wire nand_4_cse;
  wire and_84_cse;
  wire mux_14_cse;
  wire for_1_unequal_itm;
  wire and_dcpl_103;
  wire and_dcpl_109;
  wire and_dcpl_113;
  wire and_dcpl_116;
  wire and_dcpl_118;
  wire and_dcpl_121;
  wire [4:0] z_out_3;
  wire [4:0] z_out_6;
  wire [5:0] nl_z_out_6;
  wire [4:0] pntr_buf_2;
  wire [5:0] nl_pntr_buf_2;
  wire or_21_cse;
  wire for_1_for_1_for_1_for_1_nor_4_cse;
  wire or_100_cse;
  wire operator_5_false_1_acc_4_itm_5_1;
  wire operator_5_false_1_acc_3_itm_5_1;
  wire operator_5_false_1_acc_2_itm_5_1;
  wire operator_5_false_1_acc_1_itm_5_1;
  wire operator_5_false_1_acc_itm_5_1;
  wire mux_53_cse;
  wire mux_54_cse;

  wire[4:0] tile_bound_mux1h_4_nl;
  wire[4:0] for_2_if_acc_nl;
  wire[5:0] nl_for_2_if_acc_nl;
  wire[4:0] for_2_if_mux_6_nl;
  wire[0:0] tile_bound_or_nl;
  wire[4:0] tile_bound_mux1h_3_nl;
  wire[4:0] for_2_if_for_acc_nl;
  wire[5:0] nl_for_2_if_for_acc_nl;
  wire[4:0] for_2_if_for_for_2_if_for_mux_5_nl;
  wire[0:0] and_175_nl;
  wire[0:0] tile_bound_or_1_nl;
  wire[4:0] tile_bound_mux1h_2_nl;
  wire[4:0] acc_nl;
  wire[5:0] nl_acc_nl;
  wire[4:0] for_2_if_for_for_2_if_for_mux_7_nl;
  wire[0:0] and_177_nl;
  wire[0:0] tile_bound_or_2_nl;
  wire[4:0] tile_bound_mux1h_1_nl;
  wire[4:0] for_2_if_for_acc_12_nl;
  wire[5:0] nl_for_2_if_for_acc_12_nl;
  wire[4:0] for_2_if_for_for_2_if_for_mux_6_nl;
  wire[0:0] and_176_nl;
  wire[0:0] tile_bound_or_3_nl;
  wire[4:0] tile_bound_mux1h_nl;
  wire[4:0] for_2_if_for_acc_13_nl;
  wire[5:0] nl_for_2_if_for_acc_13_nl;
  wire[4:0] for_2_if_for_for_2_if_for_mux_4_nl;
  wire[0:0] and_174_nl;
  wire[0:0] mux_52_nl;
  wire[0:0] tile_bound_or_4_nl;
  wire[4:0] tile_pntr_and_nl;
  wire[0:0] tile_pntr_nand_nl;
  wire[0:0] mux_44_nl;
  wire[0:0] mux_43_nl;
  wire[0:0] mux_42_nl;
  wire[0:0] mux_41_nl;
  wire[0:0] mux_40_nl;
  wire[0:0] mux_39_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] and_88_nl;
  wire[4:0] for_2_if_for_for_2_if_for_and_1_nl;
  wire[4:0] for_2_if_for_mux_1_nl;
  wire[0:0] nor_24_nl;
  wire[0:0] counter_nand_4_nl;
  wire[0:0] mux_24_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] nor_21_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] mux_21_nl;
  wire[0:0] nand_3_nl;
  wire[0:0] or_26_nl;
  wire[0:0] or_24_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] mux_32_nl;
  wire[0:0] mux_31_nl;
  wire[0:0] nor_18_nl;
  wire[0:0] mux_30_nl;
  wire[0:0] nand_1_nl;
  wire[0:0] or_44_nl;
  wire[0:0] mux_29_nl;
  wire[0:0] nor_5_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] mux_37_nl;
  wire[0:0] mux_36_nl;
  wire[0:0] or_59_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] or_56_nl;
  wire[0:0] mux_34_nl;
  wire[0:0] nor_7_nl;
  wire[0:0] mux_45_nl;
  wire[0:0] nor_30_nl;
  wire[0:0] nand_7_nl;
  wire[0:0] nor_10_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] mux_10_nl;
  wire[4:0] for_2_if_for_mux_nl;
  wire[0:0] counter_nand_3_nl;
  wire[4:0] for_2_if_for_mux_2_nl;
  wire[0:0] counter_nand_2_nl;
  wire[4:0] for_2_if_for_mux_3_nl;
  wire[0:0] counter_nand_1_nl;
  wire[4:0] for_2_if_for_mux_4_nl;
  wire[0:0] counter_or_nl;
  wire[4:0] counter_mux_nl;
  wire[0:0] counter_nand_nl;
  wire[5:0] operator_5_false_1_acc_4_nl;
  wire[6:0] nl_operator_5_false_1_acc_4_nl;
  wire[5:0] operator_5_false_1_acc_3_nl;
  wire[6:0] nl_operator_5_false_1_acc_3_nl;
  wire[5:0] operator_5_false_1_acc_2_nl;
  wire[6:0] nl_operator_5_false_1_acc_2_nl;
  wire[5:0] operator_5_false_1_acc_1_nl;
  wire[6:0] nl_operator_5_false_1_acc_1_nl;
  wire[5:0] operator_5_false_1_acc_nl;
  wire[6:0] nl_operator_5_false_1_acc_nl;
  wire[0:0] nand_nl;
  wire[0:0] or_34_nl;
  wire[0:0] mux_26_nl;
  wire[0:0] mux_25_nl;
  wire[0:0] or_32_nl;
  wire[0:0] or_31_nl;
  wire[0:0] and_171_nl;
  wire[5:0] acc_3_nl;
  wire[6:0] nl_acc_3_nl;
  wire[4:0] for_2_if_mux1h_3_nl;
  wire[4:0] for_2_if_mux1h_4_nl;
  wire[4:0] for_2_if_mux1h_5_nl;
  wire[0:0] and_179_nl;

  // Interconnect Declarations for Component Instantiations 
  assign counter_out = {counter_buf_4_1_mx0 , counter_buf_3_1_mx0 , counter_buf_2_1_mx0
      , counter_buf_1_1_mx0 , counter_buf_0_1_mx1};
  assign for_2_if_mux_6_nl = MUX_v_5_2_2(z_out_3, (tile_bound_in[24:20]), for_1_for_1_for_1_for_1_nor_4_cse);
  assign nl_for_2_if_acc_nl = for_2_if_mux_6_nl + (tile_sizes[24:20]);
  assign for_2_if_acc_nl = nl_for_2_if_acc_nl[4:0];
  assign tile_bound_or_nl = and_dcpl_53 | (and_dcpl_64 & (~ equal_mdf_1) & operator_5_false_1_acc_4_itm_5_1
      & (~ for_1_unequal_3_tmp) & and_dcpl);
  assign tile_bound_mux1h_4_nl = MUX1HOT_v_5_3_2(for_2_if_acc_nl, (tile_sizes[24:20]),
      (tile_bound_in[24:20]), {tile_bound_or_nl , and_dcpl_65 , or_dcpl_25});
  assign and_175_nl = (~(or_82_cse & operator_5_false_1_acc_4_itm_5_1)) & and_dcpl_103;
  assign for_2_if_for_for_2_if_for_mux_5_nl = MUX_v_5_2_2(z_out_3, (tile_bound_in[19:15]),
      and_175_nl);
  assign nl_for_2_if_for_acc_nl = for_2_if_for_for_2_if_for_mux_5_nl + (tile_sizes[19:15]);
  assign for_2_if_for_acc_nl = nl_for_2_if_for_acc_nl[4:0];
  assign tile_bound_or_1_nl = and_dcpl_53 | and_dcpl_46 | ((nor_16_cse | (~ operator_5_false_1_acc_4_itm_5_1))
      & and_dcpl_3 & and_dcpl_12 & operator_5_false_1_acc_3_itm_5_1 & and_dcpl_38);
  assign tile_bound_mux1h_3_nl = MUX1HOT_v_5_3_2(for_2_if_for_acc_nl, (tile_sizes[19:15]),
      (tile_bound_in[19:15]), {tile_bound_or_1_nl , and_dcpl_65 , or_dcpl_21});
  assign and_177_nl = (~ mux_54_cse) & and_dcpl_12;
  assign for_2_if_for_for_2_if_for_mux_7_nl = MUX_v_5_2_2(z_out_3, (tile_bound_in[14:10]),
      and_177_nl);
  assign nl_acc_nl = for_2_if_for_for_2_if_for_mux_7_nl + (tile_sizes[14:10]);
  assign acc_nl = nl_acc_nl[4:0];
  assign tile_bound_or_2_nl = and_dcpl_53 | and_dcpl_46 | and_dcpl_35 | ((~ mux_tmp_30)
      & and_dcpl_4 & (~ (operator_5_false_acc_2_tmp[5])) & operator_5_false_1_acc_2_itm_5_1
      & for_1_for_1_for_1_for_1_nor_tmp);
  assign tile_bound_mux1h_2_nl = MUX1HOT_v_5_3_2(acc_nl, (tile_sizes[14:10]), (tile_bound_in[14:10]),
      {tile_bound_or_2_nl , and_dcpl_65 , or_dcpl_13});
  assign and_176_nl = (~ mux_53_cse) & and_dcpl_3;
  assign for_2_if_for_for_2_if_for_mux_6_nl = MUX_v_5_2_2(z_out_3, (tile_bound_in[9:5]),
      and_176_nl);
  assign nl_for_2_if_for_acc_12_nl = for_2_if_for_for_2_if_for_mux_6_nl + (tile_sizes[9:5]);
  assign for_2_if_for_acc_12_nl = nl_for_2_if_for_acc_12_nl[4:0];
  assign tile_bound_or_3_nl = and_dcpl_53 | and_dcpl_46 | and_dcpl_35 | and_dcpl_28
      | ((~ mux_tmp_25) & and_dcpl_3 & and_dcpl_27);
  assign tile_bound_mux1h_1_nl = MUX1HOT_v_5_3_2(for_2_if_for_acc_12_nl, (tile_sizes[9:5]),
      (tile_bound_in[9:5]), {tile_bound_or_3_nl , and_dcpl_65 , or_dcpl_10});
  assign mux_52_nl = MUX_s_1_2_2(mux_53_cse, operator_5_false_1_acc_1_itm_5_1, or_20_cse);
  assign and_174_nl = (~ mux_52_nl) & for_1_for_1_for_1_for_1_nor_tmp;
  assign for_2_if_for_for_2_if_for_mux_4_nl = MUX_v_5_2_2(z_out_3, (tile_bound_in[4:0]),
      and_174_nl);
  assign nl_for_2_if_for_acc_13_nl = for_2_if_for_for_2_if_for_mux_4_nl + (tile_sizes[4:0]);
  assign for_2_if_for_acc_13_nl = nl_for_2_if_for_acc_13_nl[4:0];
  assign tile_bound_or_4_nl = and_dcpl_53 | and_dcpl_46 | and_dcpl_35 | and_dcpl_28
      | ((~ for_1_for_1_for_1_for_1_nor_tmp) & operator_5_false_1_acc_itm_5_1) |
      ((~ mux_14_cse) & for_1_for_1_for_1_for_1_nor_tmp & operator_5_false_1_acc_itm_5_1);
  assign tile_bound_mux1h_nl = MUX1HOT_v_5_3_2(for_2_if_for_acc_13_nl, (tile_sizes[4:0]),
      (tile_bound_in[4:0]), {tile_bound_or_4_nl , and_dcpl_65 , and_dcpl_24});
  assign tile_bound_out = {tile_bound_mux1h_4_nl , tile_bound_mux1h_3_nl , tile_bound_mux1h_2_nl
      , tile_bound_mux1h_1_nl , tile_bound_mux1h_nl};
  assign or_89_cse = equal_mdf_1 | for_1_unequal_4_tmp | (operator_5_false_acc_4_tmp[5]);
  assign or_79_cse = for_1_unequal_3_tmp | (operator_5_false_acc_3_tmp[5]);
  assign or_75_cse = for_1_unequal_2_tmp | (operator_5_false_acc_2_tmp[5]);
  assign and_84_cse = or_89_cse & operator_5_false_1_acc_4_itm_5_1;
  assign tile_pntr_nand_nl = ~(and_dcpl_10 & (~ (operator_5_false_acc_4_tmp[5]))
      & (~ for_1_unequal_3_tmp) & and_dcpl);
  assign tile_pntr_and_nl = MUX_v_5_2_2(5'b00000, z_out_3, tile_pntr_nand_nl);
  assign mux_41_nl = MUX_s_1_2_2(and_tmp, or_tmp_48, and_84_cse);
  assign mux_40_nl = MUX_s_1_2_2(and_tmp, or_tmp_48, operator_5_false_1_acc_3_itm_5_1);
  assign mux_42_nl = MUX_s_1_2_2(mux_41_nl, mux_40_nl, or_79_cse);
  assign mux_39_nl = MUX_s_1_2_2(and_tmp, or_tmp_48, operator_5_false_1_acc_2_itm_5_1);
  assign mux_43_nl = MUX_s_1_2_2(mux_42_nl, mux_39_nl, or_75_cse);
  assign mux_44_nl = MUX_s_1_2_2(operator_5_false_1_acc_itm_5_1, mux_43_nl, for_1_for_1_for_1_for_1_nor_tmp);
  assign pntr_out = MUX_v_5_2_2(pntr_buf_2, tile_pntr_and_nl, mux_44_nl);
  assign and_88_nl = (equal_mdf_1 | for_1_unequal_4_tmp) & operator_5_false_1_acc_4_itm_5_1;
  assign mux_7_nl = MUX_s_1_2_2(and_88_nl, operator_5_false_1_acc_3_itm_5_1, for_1_unequal_3_tmp);
  assign mux_8_nl = MUX_s_1_2_2(mux_7_nl, operator_5_false_1_acc_2_itm_5_1, for_1_unequal_2_tmp);
  assign mux_9_cse = MUX_s_1_2_2(mux_8_nl, operator_5_false_1_acc_1_itm_5_1, for_1_unequal_1_tmp);
  assign nor_24_nl = ~((mux_9_cse & for_1_for_1_for_1_for_1_nor_tmp) | operator_5_false_1_acc_itm_5_1);
  assign for_2_if_for_mux_1_nl = MUX_v_5_2_2(z_out_6, (counter_in[4:0]), nor_24_nl);
  assign counter_nand_4_nl = ~((mux_9_cse | operator_5_false_1_acc_itm_5_1) & for_1_for_1_for_1_for_1_nor_tmp);
  assign for_2_if_for_for_2_if_for_and_1_nl = MUX_v_5_2_2(5'b00000, for_2_if_for_mux_1_nl,
      counter_nand_4_nl);
  assign irrel_at_max_out = (~((for_2_if_for_for_2_if_for_and_1_nl != (operator_5_false_acc_cse_1[4:0]))
      | (operator_5_false_acc_cse_1[5]))) & (~((operator_5_false_acc_1_tmp[5]) |
      (counter_buf_1_1_mx0 != (operator_5_false_acc_1_tmp[4:0])))) & (~((operator_5_false_acc_2_tmp[5])
      | (counter_buf_2_1_mx0 != (operator_5_false_acc_2_tmp[4:0])))) & (~((operator_5_false_acc_3_tmp[5])
      | (counter_buf_3_1_mx0 != (operator_5_false_acc_3_tmp[4:0])))) & (~((operator_5_false_acc_4_tmp[5])
      | (counter_buf_4_1_mx0 != (operator_5_false_acc_4_tmp[4:0]))));
  assign or_82_cse = for_1_unequal_4_tmp | (operator_5_false_acc_4_tmp[5]);
  assign or_20_cse = for_1_unequal_1_tmp | (operator_5_false_acc_1_tmp[5]);
  assign nor_16_cse = ~(equal_mdf_1 | for_1_unequal_4_tmp | (operator_5_false_acc_4_tmp[5]));
  assign nand_4_cse = ~(or_89_cse & operator_5_false_1_acc_4_itm_5_1);
  assign or_21_cse = (z_out_6!=5'b00000);
  assign nand_3_nl = ~(nand_4_cse & or_tmp_14);
  assign or_26_nl = operator_5_false_1_acc_3_itm_5_1 | (~ or_tmp_14);
  assign mux_21_nl = MUX_s_1_2_2(nand_3_nl, or_26_nl, or_79_cse);
  assign or_24_nl = operator_5_false_1_acc_2_itm_5_1 | (~ or_tmp_14);
  assign mux_22_nl = MUX_s_1_2_2(mux_21_nl, or_24_nl, or_75_cse);
  assign nor_21_nl = ~(operator_5_false_1_acc_1_itm_5_1 | mux_22_nl);
  assign mux_20_nl = MUX_s_1_2_2(or_tmp_14, or_21_cse, operator_5_false_1_acc_1_itm_5_1);
  assign mux_23_nl = MUX_s_1_2_2(nor_21_nl, mux_20_nl, or_20_cse);
  assign mux_24_nl = MUX_s_1_2_2(or_tmp_14, mux_23_nl, for_1_for_1_for_1_for_1_nor_tmp);
  assign nand_1_nl = ~(nand_4_cse & or_tmp_31);
  assign or_44_nl = operator_5_false_1_acc_3_itm_5_1 | (~ or_tmp_31);
  assign mux_30_nl = MUX_s_1_2_2(nand_1_nl, or_44_nl, or_79_cse);
  assign nor_18_nl = ~(operator_5_false_1_acc_2_itm_5_1 | mux_30_nl);
  assign mux_29_nl = MUX_s_1_2_2(or_tmp_31, or_21_cse, operator_5_false_1_acc_2_itm_5_1);
  assign mux_31_nl = MUX_s_1_2_2(nor_18_nl, mux_29_nl, or_75_cse);
  assign nor_5_nl = ~(for_1_unequal_1_tmp | (operator_5_false_acc_1_tmp[5]) | (~
      for_1_for_1_for_1_for_1_nor_tmp));
  assign mux_32_nl = MUX_s_1_2_2(or_tmp_31, mux_31_nl, nor_5_nl);
  assign or_59_nl = nor_16_cse | (~ operator_5_false_1_acc_4_itm_5_1) | for_1_unequal_2_tmp
      | (operator_5_false_acc_2_tmp[5]) | for_1_unequal_1_tmp | (operator_5_false_acc_1_tmp[5]);
  assign mux_36_nl = MUX_s_1_2_2(not_tmp_24, or_tmp_41, or_59_nl);
  assign or_56_nl = for_1_unequal_2_tmp | (operator_5_false_acc_2_tmp[5]) | for_1_unequal_1_tmp
      | (operator_5_false_acc_1_tmp[5]);
  assign mux_35_nl = MUX_s_1_2_2(not_tmp_24, or_tmp_41, or_56_nl);
  assign mux_37_nl = MUX_s_1_2_2(mux_36_nl, mux_35_nl, operator_5_false_1_acc_3_itm_5_1);
  assign nor_7_nl = ~((~ operator_5_false_1_acc_3_itm_5_1) | for_1_unequal_2_tmp
      | (operator_5_false_acc_2_tmp[5]) | for_1_unequal_1_tmp | (operator_5_false_acc_1_tmp[5])
      | (~ for_1_for_1_for_1_for_1_nor_tmp));
  assign mux_34_nl = MUX_s_1_2_2(or_tmp_41, or_21_cse, nor_7_nl);
  assign mux_38_nl = MUX_s_1_2_2(mux_37_nl, mux_34_nl, or_79_cse);
  assign nor_30_nl = ~((counter_in[24:20]!=5'b00000));
  assign nand_7_nl = ~(or_82_cse & or_21_cse);
  assign nor_10_nl = ~((~ operator_5_false_1_acc_4_itm_5_1) | for_1_unequal_3_tmp
      | (operator_5_false_acc_3_tmp[5]) | for_1_unequal_2_tmp | (operator_5_false_acc_2_tmp[5])
      | for_1_unequal_1_tmp | (operator_5_false_acc_1_tmp[5]) | (~ for_1_for_1_for_1_for_1_nor_tmp));
  assign mux_45_nl = MUX_s_1_2_2(nor_30_nl, nand_7_nl, nor_10_nl);
  assign irrel_at_zero_out = (~((counter_buf_0_1_mx1!=5'b00000) | mux_24_nl | mux_32_nl
      | mux_38_nl)) & mux_45_nl;
  assign for_1_for_1_for_1_for_1_nor_4_cse = ~(for_1_unequal_4_tmp | (operator_5_false_acc_4_tmp[5]));
  assign all_at_max_1_out = for_1_for_1_for_1_for_1_nor_4_cse & (~(or_dcpl_16 | (operator_5_false_acc_2_tmp[5])
      | (~ equal_mdf_1) | or_dcpl_23));
  assign mux_12_nl = MUX_s_1_2_2(and_tmp, or_tmp_4, and_84_cse);
  assign mux_11_nl = MUX_s_1_2_2(and_tmp, or_tmp_4, operator_5_false_1_acc_3_itm_5_1);
  assign mux_13_nl = MUX_s_1_2_2(mux_12_nl, mux_11_nl, or_79_cse);
  assign mux_10_nl = MUX_s_1_2_2(and_tmp, or_tmp_4, operator_5_false_1_acc_2_itm_5_1);
  assign mux_14_cse = MUX_s_1_2_2(mux_13_nl, mux_10_nl, or_75_cse);
  assign for_2_if_for_mux_nl = MUX_v_5_2_2(z_out_6, (counter_in[4:0]), and_dcpl_24);
  assign counter_nand_3_nl = ~((mux_14_cse | operator_5_false_1_acc_itm_5_1) & for_1_for_1_for_1_for_1_nor_tmp);
  assign counter_buf_0_1_mx1 = MUX_v_5_2_2(5'b00000, for_2_if_for_mux_nl, counter_nand_3_nl);
  assign for_2_if_for_mux_2_nl = MUX_v_5_2_2(z_out_6, (counter_in[9:5]), or_dcpl_10);
  assign counter_nand_2_nl = ~((mux_tmp_25 | operator_5_false_1_acc_1_itm_5_1) &
      and_dcpl_3 & for_1_for_1_for_1_for_1_nor_tmp);
  assign counter_buf_1_1_mx0 = MUX_v_5_2_2(5'b00000, for_2_if_for_mux_2_nl, counter_nand_2_nl);
  assign nl_pntr_buf_2 = pntr_in + 5'b00001;
  assign pntr_buf_2 = nl_pntr_buf_2[4:0];
  assign for_2_if_for_mux_3_nl = MUX_v_5_2_2(z_out_6, (counter_in[14:10]), or_dcpl_13);
  assign counter_nand_1_nl = ~((mux_tmp_30 | operator_5_false_1_acc_2_itm_5_1) &
      and_dcpl_4 & (~ (operator_5_false_acc_2_tmp[5])) & for_1_for_1_for_1_for_1_nor_tmp);
  assign counter_buf_2_1_mx0 = MUX_v_5_2_2(5'b00000, for_2_if_for_mux_3_nl, counter_nand_1_nl);
  assign for_2_if_for_mux_4_nl = MUX_v_5_2_2(z_out_6, (counter_in[19:15]), or_dcpl_21);
  assign counter_or_nl = (~(and_84_cse | operator_5_false_1_acc_3_itm_5_1)) | for_1_unequal_1_tmp
      | (operator_5_false_acc_1_tmp[5]) | for_1_unequal_2_tmp | (operator_5_false_acc_2_tmp[5])
      | (~ and_dcpl_38);
  assign counter_buf_3_1_mx0 = MUX_v_5_2_2(5'b00000, for_2_if_for_mux_4_nl, counter_or_nl);
  assign counter_mux_nl = MUX_v_5_2_2(z_out_6, (counter_in[24:20]), or_dcpl_25);
  assign counter_nand_nl = ~(and_dcpl_10 & (~ (operator_5_false_acc_4_tmp[5])) &
      operator_5_false_1_acc_4_itm_5_1 & (~ for_1_unequal_3_tmp) & and_dcpl);
  assign counter_buf_4_1_mx0 = MUX_v_5_2_2(5'b00000, counter_mux_nl, counter_nand_nl);
  assign for_1_unequal_4_tmp = (counter_in[24:20]) != (operator_5_false_acc_4_tmp[4:0]);
  assign nl_operator_5_false_acc_cse_1 = conv_u2s_5_6(loop_bound[4:0]) + 6'b111111;
  assign operator_5_false_acc_cse_1 = nl_operator_5_false_acc_cse_1[5:0];
  assign nl_operator_5_false_acc_4_tmp = conv_u2s_5_6(loop_bound[24:20]) + 6'b111111;
  assign operator_5_false_acc_4_tmp = nl_operator_5_false_acc_4_tmp[5:0];
  assign nl_operator_5_false_acc_3_tmp = conv_u2s_5_6(loop_bound[19:15]) + 6'b111111;
  assign operator_5_false_acc_3_tmp = nl_operator_5_false_acc_3_tmp[5:0];
  assign nl_operator_5_false_acc_2_tmp = conv_u2s_5_6(loop_bound[14:10]) + 6'b111111;
  assign operator_5_false_acc_2_tmp = nl_operator_5_false_acc_2_tmp[5:0];
  assign nl_operator_5_false_acc_1_tmp = conv_u2s_5_6(loop_bound[9:5]) + 6'b111111;
  assign operator_5_false_acc_1_tmp = nl_operator_5_false_acc_1_tmp[5:0];
  assign equal_mdf_1 = pntr_buf_2 == (tile_sizes[24:20]);
  assign nl_operator_5_false_1_acc_4_nl = ({1'b1 , (tile_bound_in[24:20])}) + conv_u2s_5_6(~
      pntr_buf_2);
  assign operator_5_false_1_acc_4_nl = nl_operator_5_false_1_acc_4_nl[5:0];
  assign operator_5_false_1_acc_4_itm_5_1 = readslicef_6_1_5(operator_5_false_1_acc_4_nl);
  assign nl_operator_5_false_1_acc_3_nl = ({1'b1 , (tile_bound_in[19:15])}) + conv_u2s_5_6(~
      pntr_buf_2);
  assign operator_5_false_1_acc_3_nl = nl_operator_5_false_1_acc_3_nl[5:0];
  assign operator_5_false_1_acc_3_itm_5_1 = readslicef_6_1_5(operator_5_false_1_acc_3_nl);
  assign for_1_unequal_3_tmp = (counter_in[19:15]) != (operator_5_false_acc_3_tmp[4:0]);
  assign nl_operator_5_false_1_acc_2_nl = ({1'b1 , (tile_bound_in[14:10])}) + conv_u2s_5_6(~
      pntr_buf_2);
  assign operator_5_false_1_acc_2_nl = nl_operator_5_false_1_acc_2_nl[5:0];
  assign operator_5_false_1_acc_2_itm_5_1 = readslicef_6_1_5(operator_5_false_1_acc_2_nl);
  assign for_1_unequal_2_tmp = (counter_in[14:10]) != (operator_5_false_acc_2_tmp[4:0]);
  assign nl_operator_5_false_1_acc_1_nl = ({1'b1 , (tile_bound_in[9:5])}) + conv_u2s_5_6(~
      pntr_buf_2);
  assign operator_5_false_1_acc_1_nl = nl_operator_5_false_1_acc_1_nl[5:0];
  assign operator_5_false_1_acc_1_itm_5_1 = readslicef_6_1_5(operator_5_false_1_acc_1_nl);
  assign for_1_unequal_1_tmp = (counter_in[9:5]) != (operator_5_false_acc_1_tmp[4:0]);
  assign nl_operator_5_false_1_acc_nl = ({1'b1 , (tile_bound_in[4:0])}) + conv_u2s_5_6(~
      pntr_buf_2);
  assign operator_5_false_1_acc_nl = nl_operator_5_false_1_acc_nl[5:0];
  assign operator_5_false_1_acc_itm_5_1 = readslicef_6_1_5(operator_5_false_1_acc_nl);
  assign for_1_unequal_itm = (counter_in[4:0]) != (operator_5_false_acc_cse_1[4:0]);
  assign for_1_for_1_for_1_for_1_nor_tmp = ~(for_1_unequal_itm | (operator_5_false_acc_cse_1[5]));
  assign and_dcpl = (~ (operator_5_false_acc_3_tmp[5])) & for_1_for_1_for_1_for_1_nor_tmp;
  assign and_dcpl_3 = ~(for_1_unequal_1_tmp | (operator_5_false_acc_1_tmp[5]));
  assign and_dcpl_4 = and_dcpl_3 & (~ for_1_unequal_2_tmp);
  assign and_dcpl_9 = ~((operator_5_false_acc_2_tmp[5]) | for_1_unequal_4_tmp);
  assign and_dcpl_10 = and_dcpl_4 & and_dcpl_9;
  assign and_dcpl_12 = ~(for_1_unequal_2_tmp | (operator_5_false_acc_2_tmp[5]));
  assign or_tmp_4 = operator_5_false_1_acc_1_itm_5_1 | (~ or_20_cse);
  assign and_tmp = operator_5_false_1_acc_1_itm_5_1 & or_20_cse;
  assign and_dcpl_24 = ~((mux_14_cse & for_1_for_1_for_1_for_1_nor_tmp) | operator_5_false_1_acc_itm_5_1);
  assign or_tmp_14 = (counter_in[9:5]!=5'b00000);
  assign nand_nl = ~(operator_5_false_1_acc_4_itm_5_1 & (~(nor_16_cse | (operator_5_false_acc_2_tmp[5])
      | for_1_unequal_2_tmp)));
  assign or_34_nl = (~ operator_5_false_1_acc_3_itm_5_1) | (operator_5_false_acc_2_tmp[5])
      | for_1_unequal_2_tmp;
  assign mux_tmp_24 = MUX_s_1_2_2(nand_nl, or_34_nl, or_79_cse);
  assign or_32_nl = equal_mdf_1 | (operator_5_false_acc_4_tmp[5]) | for_1_unequal_4_tmp
      | (operator_5_false_acc_2_tmp[5]) | for_1_unequal_2_tmp;
  assign mux_25_nl = MUX_s_1_2_2(or_75_cse, or_32_nl, operator_5_false_1_acc_4_itm_5_1);
  assign or_31_nl = operator_5_false_1_acc_3_itm_5_1 | (operator_5_false_acc_2_tmp[5])
      | for_1_unequal_2_tmp;
  assign mux_26_nl = MUX_s_1_2_2(mux_25_nl, or_31_nl, or_79_cse);
  assign mux_tmp_25 = MUX_s_1_2_2((~ mux_tmp_24), mux_26_nl, operator_5_false_1_acc_2_itm_5_1);
  assign and_dcpl_27 = operator_5_false_1_acc_1_itm_5_1 & for_1_for_1_for_1_for_1_nor_tmp;
  assign and_dcpl_28 = or_20_cse & and_dcpl_27;
  assign or_dcpl_10 = ~(((~((~ mux_tmp_25) | or_20_cse)) | operator_5_false_1_acc_1_itm_5_1)
      & for_1_for_1_for_1_for_1_nor_tmp);
  assign or_tmp_31 = (counter_in[14:10]!=5'b00000);
  assign mux_tmp_30 = MUX_s_1_2_2(and_84_cse, operator_5_false_1_acc_3_itm_5_1, or_79_cse);
  assign and_dcpl_35 = or_75_cse & (~ for_1_unequal_1_tmp) & (~ (operator_5_false_acc_1_tmp[5]))
      & operator_5_false_1_acc_2_itm_5_1 & for_1_for_1_for_1_for_1_nor_tmp;
  assign or_dcpl_13 = (mux_tmp_24 & (~ operator_5_false_1_acc_2_itm_5_1)) | or_20_cse
      | (~ for_1_for_1_for_1_for_1_nor_tmp);
  assign or_tmp_41 = (counter_in[19:15]!=5'b00000);
  assign not_tmp_24 = ~(for_1_for_1_for_1_for_1_nor_tmp | (~ or_tmp_41));
  assign and_dcpl_38 = (~ for_1_unequal_3_tmp) & (~ (operator_5_false_acc_3_tmp[5]))
      & for_1_for_1_for_1_for_1_nor_tmp;
  assign and_dcpl_46 = and_dcpl_3 & or_79_cse & and_dcpl_12 & operator_5_false_1_acc_3_itm_5_1
      & for_1_for_1_for_1_for_1_nor_tmp;
  assign or_dcpl_16 = or_20_cse | for_1_unequal_2_tmp;
  assign or_dcpl_18 = (~ operator_5_false_1_acc_4_itm_5_1) | for_1_unequal_3_tmp;
  assign or_dcpl_21 = (~((~(nor_16_cse | or_dcpl_18 | (operator_5_false_acc_3_tmp[5])))
      | operator_5_false_1_acc_3_itm_5_1)) | or_dcpl_16 | (operator_5_false_acc_2_tmp[5])
      | (~ for_1_for_1_for_1_for_1_nor_tmp);
  assign and_dcpl_53 = and_dcpl_4 & or_82_cse & (~ (operator_5_false_acc_2_tmp[5]))
      & operator_5_false_1_acc_4_itm_5_1 & (~ for_1_unequal_3_tmp) & and_dcpl;
  assign or_dcpl_23 = or_dcpl_18 | (operator_5_false_acc_3_tmp[5]) | (~ for_1_for_1_for_1_for_1_nor_tmp);
  assign or_dcpl_25 = or_20_cse | or_75_cse | or_dcpl_23;
  assign or_tmp_48 = and_dcpl_3 | operator_5_false_1_acc_1_itm_5_1;
  assign and_dcpl_64 = and_dcpl_4 & and_dcpl_9 & (~ (operator_5_false_acc_4_tmp[5]));
  assign and_dcpl_65 = and_dcpl_64 & equal_mdf_1 & operator_5_false_1_acc_4_itm_5_1
      & (~ for_1_unequal_3_tmp) & and_dcpl;
  assign or_100_cse = (operator_5_false_acc_cse_1[5]) | for_1_unequal_itm;
  assign and_dcpl_103 = ~((operator_5_false_acc_3_tmp[5]) | for_1_unequal_3_tmp);
  assign and_dcpl_109 = for_1_for_1_for_1_for_1_nor_tmp & or_20_cse;
  assign and_dcpl_113 = ~(and_dcpl_12 | (operator_5_false_acc_cse_1[5]) | for_1_unequal_itm
      | (operator_5_false_acc_1_tmp[5]) | for_1_unequal_1_tmp);
  assign and_dcpl_116 = ~((operator_5_false_acc_2_tmp[5]) | for_1_unequal_2_tmp |
      (operator_5_false_acc_1_tmp[5]) | for_1_unequal_1_tmp);
  assign and_dcpl_118 = for_1_for_1_for_1_for_1_nor_tmp & or_79_cse & and_dcpl_116;
  assign and_dcpl_121 = for_1_for_1_for_1_for_1_nor_tmp & and_dcpl_103 & and_dcpl_116;
  assign and_171_nl = or_82_cse & operator_5_false_1_acc_4_itm_5_1;
  assign mux_54_cse = MUX_s_1_2_2(and_171_nl, operator_5_false_1_acc_3_itm_5_1, or_79_cse);
  assign mux_53_cse = MUX_s_1_2_2(mux_54_cse, operator_5_false_1_acc_2_itm_5_1, or_75_cse);
  assign for_2_if_mux1h_3_nl = MUX1HOT_v_5_5_2((tile_bound_in[4:0]), (tile_bound_in[9:5]),
      (tile_bound_in[14:10]), (tile_bound_in[19:15]), (tile_bound_in[24:20]), {or_100_cse
      , and_dcpl_109 , and_dcpl_113 , and_dcpl_118 , and_dcpl_121});
  assign for_2_if_mux1h_4_nl = MUX1HOT_v_5_5_2((~ (tile_sizes[4:0])), (~ (tile_sizes[9:5])),
      (~ (tile_sizes[14:10])), (~ (tile_sizes[19:15])), (~ (tile_sizes[24:20])),
      {or_100_cse , and_dcpl_109 , and_dcpl_113 , and_dcpl_118 , and_dcpl_121});
  assign nl_acc_3_nl = ({for_2_if_mux1h_3_nl , 1'b1}) + ({for_2_if_mux1h_4_nl , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[5:0];
  assign z_out_3 = readslicef_6_5_1(acc_3_nl);
  assign and_179_nl = (~(and_dcpl_12 | for_1_unequal_itm)) & (~((operator_5_false_acc_cse_1[5])
      | (operator_5_false_acc_1_tmp[5]) | for_1_unequal_1_tmp));
  assign for_2_if_mux1h_5_nl = MUX1HOT_v_5_5_2((counter_in[4:0]), (counter_in[9:5]),
      (counter_in[14:10]), (counter_in[19:15]), (counter_in[24:20]), {or_100_cse
      , and_dcpl_109 , and_179_nl , and_dcpl_118 , and_dcpl_121});
  assign nl_z_out_6 = for_2_if_mux1h_5_nl + 5'b00001;
  assign z_out_6 = nl_z_out_6[4:0];

  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_5_2;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [4:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    result = result | ( input_3 & {5{sel[3]}});
    result = result | ( input_4 & {5{sel[4]}});
    MUX1HOT_v_5_5_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function automatic [4:0] readslicef_6_5_1;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_6_5_1 = tmp[4:0];
  end
  endfunction


  function automatic [5:0] conv_u2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_6 =  {1'b0, vector};
  end
  endfunction

endmodule




//------> /esat/micas-data/software/Mentor/catapult_10.5c/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /esat/micas-data/software/Mentor/catapult_10.5c/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ../td_ccore_solutions/tiling_unit_5_W_addr_type_L3__70f247a0b6d72f8412d9d2d7bfe58aa0b849_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   r0678912@amazone.esat.kuleuven.be
//  Generated date: Tue Jul 13 10:57:37 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    tiling_unit_5_W_addr_type_L3_run
// ------------------------------------------------------------------


module tiling_unit_5_W_addr_type_L3_run (
  loops_bound_rsc_dat, loops_relevancy_rsc_dat, tile_size_in_rsc_dat, tile_size_out_rsc_z,
      instr_bound_rsc_z, instr_tile_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [79:0] loops_bound_rsc_dat;
  input [4:0] loops_relevancy_rsc_dat;
  input [15:0] tile_size_in_rsc_dat;
  output [15:0] tile_size_out_rsc_z;
  output [79:0] instr_bound_rsc_z;
  output [79:0] instr_tile_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [79:0] loops_bound_rsci_idat;
  wire [4:0] loops_relevancy_rsci_idat;
  wire [15:0] tile_size_in_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [15:0] instr_bound_rsci_d_79_64;
  reg [15:0] instr_bound_rsci_d_63_48;
  reg [15:0] instr_bound_rsci_d_47_32;
  reg [15:0] instr_bound_rsci_d_31_16;
  reg [15:0] instr_bound_rsci_d_15_0;
  reg [4:0] instr_tile_rsci_d_15_11;
  reg [10:0] instr_tile_rsci_d_10_0;
  reg [4:0] instr_tile_rsci_d_63_59;
  reg [10:0] instr_tile_rsci_d_58_48;
  reg [4:0] instr_tile_rsci_d_47_43;
  reg [10:0] instr_tile_rsci_d_42_32;
  reg [4:0] instr_tile_rsci_d_31_27;
  reg [10:0] instr_tile_rsci_d_26_16;
  reg [4:0] reg_tile_size_out_rsci_d_15_11_cse;
  reg [10:0] reg_tile_size_out_rsci_d_10_0_cse;
  wire [10:0] instr_tile_rsci_d_10_0_mx0;
  wire [4:0] instr_tile_rsci_d_63_59_mx0;
  wire [10:0] instr_tile_rsci_d_58_48_mx0;
  wire [4:0] tile_size_int_lpi_1_dfm_15_11_1;
  wire [4:0] instr_tile_rsci_d_47_43_mx0;
  wire [10:0] instr_tile_rsci_d_42_32_mx0;
  wire [4:0] instr_tile_rsci_d_31_27_mx0;
  wire [10:0] instr_tile_rsci_d_26_16_mx0;
  wire [15:0] tile_size_int_sva_6;
  wire [26:0] nl_tile_size_int_sva_6;
  wire [15:0] tile_size_int_sva_7;
  wire [31:0] nl_tile_size_int_sva_7;
  wire [15:0] tile_size_int_sva_8;
  wire [31:0] nl_tile_size_int_sva_8;
  wire [15:0] tile_size_int_sva_9;
  wire [31:0] nl_tile_size_int_sva_9;
  wire [15:0] tile_size_int_sva_10;
  wire [31:0] nl_tile_size_int_sva_10;
  wire tile_size_and_cse;


  // Interconnect Declarations for Component Instantiations 
  wire [79:0] nl_instr_bound_rsci_d;
  assign nl_instr_bound_rsci_d = {instr_bound_rsci_d_79_64 , instr_bound_rsci_d_63_48
      , instr_bound_rsci_d_47_32 , instr_bound_rsci_d_31_16 , instr_bound_rsci_d_15_0};
  wire [79:0] nl_instr_tile_rsci_d;
  assign nl_instr_tile_rsci_d = {reg_tile_size_out_rsci_d_15_11_cse , reg_tile_size_out_rsci_d_10_0_cse
      , instr_tile_rsci_d_63_59 , instr_tile_rsci_d_58_48 , instr_tile_rsci_d_47_43
      , instr_tile_rsci_d_42_32 , instr_tile_rsci_d_31_27 , instr_tile_rsci_d_26_16
      , instr_tile_rsci_d_15_11 , instr_tile_rsci_d_10_0};
  wire [15:0] nl_tile_size_out_rsci_d;
  assign nl_tile_size_out_rsci_d = {reg_tile_size_out_rsci_d_15_11_cse , reg_tile_size_out_rsci_d_10_0_cse};
  ccs_in_v1 #(.rscid(32'sd21),
  .width(32'sd80)) loops_bound_rsci (
      .dat(loops_bound_rsc_dat),
      .idat(loops_bound_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd22),
  .width(32'sd5)) loops_relevancy_rsci (
      .dat(loops_relevancy_rsc_dat),
      .idat(loops_relevancy_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd24),
  .width(32'sd80)) instr_bound_rsci (
      .d(nl_instr_bound_rsci_d[79:0]),
      .z(instr_bound_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd25),
  .width(32'sd80)) instr_tile_rsci (
      .d(nl_instr_tile_rsci_d[79:0]),
      .z(instr_tile_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd122),
  .width(32'sd16)) tile_size_in_rsci (
      .dat(tile_size_in_rsc_dat),
      .idat(tile_size_in_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd123),
  .width(32'sd16)) tile_size_out_rsci (
      .d(nl_tile_size_out_rsci_d[15:0]),
      .z(tile_size_out_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd133),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign tile_size_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  assign instr_tile_rsci_d_10_0_mx0 = MUX_v_11_2_2((tile_size_in_rsci_idat[10:0]),
      (tile_size_int_sva_6[10:0]), loops_relevancy_rsci_idat[0]);
  assign instr_tile_rsci_d_63_59_mx0 = MUX_v_5_2_2(instr_tile_rsci_d_47_43_mx0, (tile_size_int_sva_9[15:11]),
      loops_relevancy_rsci_idat[3]);
  assign instr_tile_rsci_d_58_48_mx0 = MUX_v_11_2_2(instr_tile_rsci_d_42_32_mx0,
      (tile_size_int_sva_9[10:0]), loops_relevancy_rsci_idat[3]);
  assign tile_size_int_lpi_1_dfm_15_11_1 = MUX_v_5_2_2(5'b00000, (tile_size_int_sva_6[15:11]),
      (loops_relevancy_rsci_idat[0]));
  assign instr_tile_rsci_d_47_43_mx0 = MUX_v_5_2_2(instr_tile_rsci_d_31_27_mx0, (tile_size_int_sva_8[15:11]),
      loops_relevancy_rsci_idat[2]);
  assign instr_tile_rsci_d_42_32_mx0 = MUX_v_11_2_2(instr_tile_rsci_d_26_16_mx0,
      (tile_size_int_sva_8[10:0]), loops_relevancy_rsci_idat[2]);
  assign instr_tile_rsci_d_31_27_mx0 = MUX_v_5_2_2(tile_size_int_lpi_1_dfm_15_11_1,
      (tile_size_int_sva_7[15:11]), loops_relevancy_rsci_idat[1]);
  assign instr_tile_rsci_d_26_16_mx0 = MUX_v_11_2_2(instr_tile_rsci_d_10_0_mx0, (tile_size_int_sva_7[10:0]),
      loops_relevancy_rsci_idat[1]);
  assign nl_tile_size_int_sva_6 = (tile_size_in_rsci_idat[10:0]) * (loops_bound_rsci_idat[15:0]);
  assign tile_size_int_sva_6 = nl_tile_size_int_sva_6[15:0];
  assign nl_tile_size_int_sva_7 = ({tile_size_int_lpi_1_dfm_15_11_1 , instr_tile_rsci_d_10_0_mx0})
      * (loops_bound_rsci_idat[31:16]);
  assign tile_size_int_sva_7 = nl_tile_size_int_sva_7[15:0];
  assign nl_tile_size_int_sva_8 = ({instr_tile_rsci_d_31_27_mx0 , instr_tile_rsci_d_26_16_mx0})
      * (loops_bound_rsci_idat[47:32]);
  assign tile_size_int_sva_8 = nl_tile_size_int_sva_8[15:0];
  assign nl_tile_size_int_sva_9 = ({instr_tile_rsci_d_47_43_mx0 , instr_tile_rsci_d_42_32_mx0})
      * (loops_bound_rsci_idat[63:48]);
  assign tile_size_int_sva_9 = nl_tile_size_int_sva_9[15:0];
  assign nl_tile_size_int_sva_10 = ({instr_tile_rsci_d_63_59_mx0 , instr_tile_rsci_d_58_48_mx0})
      * (loops_bound_rsci_idat[79:64]);
  assign tile_size_int_sva_10 = nl_tile_size_int_sva_10[15:0];
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      reg_tile_size_out_rsci_d_15_11_cse <= 5'b00000;
      reg_tile_size_out_rsci_d_10_0_cse <= 11'b00000000000;
      instr_tile_rsci_d_15_11 <= 5'b00000;
    end
    else if ( tile_size_and_cse ) begin
      reg_tile_size_out_rsci_d_15_11_cse <= MUX_v_5_2_2(instr_tile_rsci_d_63_59_mx0,
          (tile_size_int_sva_10[15:11]), loops_relevancy_rsci_idat[4]);
      reg_tile_size_out_rsci_d_10_0_cse <= MUX_v_11_2_2(instr_tile_rsci_d_58_48_mx0,
          (tile_size_int_sva_10[10:0]), loops_relevancy_rsci_idat[4]);
      instr_tile_rsci_d_15_11 <= tile_size_int_lpi_1_dfm_15_11_1;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      instr_bound_rsci_d_79_64 <= 16'b0000000000000000;
      instr_bound_rsci_d_15_0 <= 16'b0000000000000000;
      instr_bound_rsci_d_63_48 <= 16'b0000000000000000;
      instr_bound_rsci_d_31_16 <= 16'b0000000000000000;
      instr_bound_rsci_d_47_32 <= 16'b0000000000000000;
      instr_tile_rsci_d_10_0 <= 11'b00000000000;
      instr_tile_rsci_d_63_59 <= 5'b00000;
      instr_tile_rsci_d_58_48 <= 11'b00000000000;
      instr_tile_rsci_d_47_43 <= 5'b00000;
      instr_tile_rsci_d_42_32 <= 11'b00000000000;
      instr_tile_rsci_d_31_27 <= 5'b00000;
      instr_tile_rsci_d_26_16 <= 11'b00000000000;
    end
    else if ( ccs_ccore_en ) begin
      instr_bound_rsci_d_79_64 <= MUX_v_16_2_2((loops_bound_rsci_idat[79:64]), 16'b0000000000000001,
          loops_relevancy_rsci_idat[4]);
      instr_bound_rsci_d_15_0 <= MUX_v_16_2_2((loops_bound_rsci_idat[15:0]), 16'b0000000000000001,
          loops_relevancy_rsci_idat[0]);
      instr_bound_rsci_d_63_48 <= MUX_v_16_2_2((loops_bound_rsci_idat[63:48]), 16'b0000000000000001,
          loops_relevancy_rsci_idat[3]);
      instr_bound_rsci_d_31_16 <= MUX_v_16_2_2((loops_bound_rsci_idat[31:16]), 16'b0000000000000001,
          loops_relevancy_rsci_idat[1]);
      instr_bound_rsci_d_47_32 <= MUX_v_16_2_2((loops_bound_rsci_idat[47:32]), 16'b0000000000000001,
          loops_relevancy_rsci_idat[2]);
      instr_tile_rsci_d_10_0 <= instr_tile_rsci_d_10_0_mx0;
      instr_tile_rsci_d_63_59 <= instr_tile_rsci_d_63_59_mx0;
      instr_tile_rsci_d_58_48 <= instr_tile_rsci_d_58_48_mx0;
      instr_tile_rsci_d_47_43 <= instr_tile_rsci_d_47_43_mx0;
      instr_tile_rsci_d_42_32 <= instr_tile_rsci_d_42_32_mx0;
      instr_tile_rsci_d_31_27 <= instr_tile_rsci_d_31_27_mx0;
      instr_tile_rsci_d_26_16 <= instr_tile_rsci_d_26_16_mx0;
    end
  end

  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    tiling_unit_5_W_addr_type_L3
// ------------------------------------------------------------------


module tiling_unit_5_W_addr_type_L3 (
  loops_bound_rsc_dat, loops_relevancy_rsc_dat, tile_size_in_rsc_dat, tile_size_out_rsc_z,
      instr_bound_rsc_z, instr_tile_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [79:0] loops_bound_rsc_dat;
  input [4:0] loops_relevancy_rsc_dat;
  input [15:0] tile_size_in_rsc_dat;
  output [15:0] tile_size_out_rsc_z;
  output [79:0] instr_bound_rsc_z;
  output [79:0] instr_tile_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  tiling_unit_5_W_addr_type_L3_run tiling_unit_5_W_addr_type_L3_run_inst (
      .loops_bound_rsc_dat(loops_bound_rsc_dat),
      .loops_relevancy_rsc_dat(loops_relevancy_rsc_dat),
      .tile_size_in_rsc_dat(tile_size_in_rsc_dat),
      .tile_size_out_rsc_z(tile_size_out_rsc_z),
      .instr_bound_rsc_z(instr_bound_rsc_z),
      .instr_tile_rsc_z(instr_tile_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/tiling_unit_5_W_addr_type_L2__207263b1b236881e25012088d06269c7b762_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   r0678912@amazone.esat.kuleuven.be
//  Generated date: Tue Jul 13 10:57:56 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    tiling_unit_5_W_addr_type_L2_run
// ------------------------------------------------------------------


module tiling_unit_5_W_addr_type_L2_run (
  loops_bound_rsc_dat, loops_relevancy_rsc_dat, tile_size_in_rsc_dat, tile_size_out_rsc_z,
      instr_bound_rsc_z, instr_tile_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [54:0] loops_bound_rsc_dat;
  input [4:0] loops_relevancy_rsc_dat;
  input [10:0] tile_size_in_rsc_dat;
  output [10:0] tile_size_out_rsc_z;
  output [54:0] instr_bound_rsc_z;
  output [54:0] instr_tile_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [54:0] loops_bound_rsci_idat;
  wire [4:0] loops_relevancy_rsci_idat;
  wire [10:0] tile_size_in_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [10:0] instr_bound_rsci_d_54_44;
  reg [10:0] instr_bound_rsci_d_43_33;
  reg [10:0] instr_bound_rsci_d_32_22;
  reg [10:0] instr_bound_rsci_d_21_11;
  reg [10:0] instr_bound_rsci_d_10_0;
  reg [5:0] instr_tile_rsci_d_10_5;
  reg [4:0] instr_tile_rsci_d_4_0;
  reg [5:0] instr_tile_rsci_d_43_38;
  reg [4:0] instr_tile_rsci_d_37_33;
  reg [5:0] instr_tile_rsci_d_32_27;
  reg [4:0] instr_tile_rsci_d_26_22;
  reg [5:0] instr_tile_rsci_d_21_16;
  reg [4:0] instr_tile_rsci_d_15_11;
  reg [5:0] reg_tile_size_out_rsci_d_10_5_cse;
  reg [4:0] reg_tile_size_out_rsci_d_4_0_cse;
  wire [4:0] instr_tile_rsci_d_4_0_mx0;
  wire [5:0] instr_tile_rsci_d_43_38_mx0;
  wire [4:0] instr_tile_rsci_d_37_33_mx0;
  wire [5:0] tile_size_int_lpi_1_dfm_10_5_1;
  wire [5:0] instr_tile_rsci_d_32_27_mx0;
  wire [4:0] instr_tile_rsci_d_26_22_mx0;
  wire [5:0] instr_tile_rsci_d_21_16_mx0;
  wire [4:0] instr_tile_rsci_d_15_11_mx0;
  wire [10:0] tile_size_int_sva_6;
  wire [15:0] nl_tile_size_int_sva_6;
  wire [10:0] tile_size_int_sva_7;
  wire [21:0] nl_tile_size_int_sva_7;
  wire [10:0] tile_size_int_sva_8;
  wire [21:0] nl_tile_size_int_sva_8;
  wire [10:0] tile_size_int_sva_9;
  wire [21:0] nl_tile_size_int_sva_9;
  wire [10:0] tile_size_int_sva_10;
  wire [21:0] nl_tile_size_int_sva_10;
  wire tile_size_and_cse;


  // Interconnect Declarations for Component Instantiations 
  wire [54:0] nl_instr_bound_rsci_d;
  assign nl_instr_bound_rsci_d = {instr_bound_rsci_d_54_44 , instr_bound_rsci_d_43_33
      , instr_bound_rsci_d_32_22 , instr_bound_rsci_d_21_11 , instr_bound_rsci_d_10_0};
  wire [54:0] nl_instr_tile_rsci_d;
  assign nl_instr_tile_rsci_d = {reg_tile_size_out_rsci_d_10_5_cse , reg_tile_size_out_rsci_d_4_0_cse
      , instr_tile_rsci_d_43_38 , instr_tile_rsci_d_37_33 , instr_tile_rsci_d_32_27
      , instr_tile_rsci_d_26_22 , instr_tile_rsci_d_21_16 , instr_tile_rsci_d_15_11
      , instr_tile_rsci_d_10_5 , instr_tile_rsci_d_4_0};
  wire [10:0] nl_tile_size_out_rsci_d;
  assign nl_tile_size_out_rsci_d = {reg_tile_size_out_rsci_d_10_5_cse , reg_tile_size_out_rsci_d_4_0_cse};
  ccs_in_v1 #(.rscid(32'sd16),
  .width(32'sd55)) loops_bound_rsci (
      .dat(loops_bound_rsc_dat),
      .idat(loops_bound_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd17),
  .width(32'sd5)) loops_relevancy_rsci (
      .dat(loops_relevancy_rsc_dat),
      .idat(loops_relevancy_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd19),
  .width(32'sd55)) instr_bound_rsci (
      .d(nl_instr_bound_rsci_d[54:0]),
      .z(instr_bound_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd20),
  .width(32'sd55)) instr_tile_rsci (
      .d(nl_instr_tile_rsci_d[54:0]),
      .z(instr_tile_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd124),
  .width(32'sd11)) tile_size_in_rsci (
      .dat(tile_size_in_rsc_dat),
      .idat(tile_size_in_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd125),
  .width(32'sd11)) tile_size_out_rsci (
      .d(nl_tile_size_out_rsci_d[10:0]),
      .z(tile_size_out_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd134),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign tile_size_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  assign instr_tile_rsci_d_4_0_mx0 = MUX_v_5_2_2((tile_size_in_rsci_idat[4:0]), (tile_size_int_sva_6[4:0]),
      loops_relevancy_rsci_idat[0]);
  assign instr_tile_rsci_d_43_38_mx0 = MUX_v_6_2_2(instr_tile_rsci_d_32_27_mx0, (tile_size_int_sva_9[10:5]),
      loops_relevancy_rsci_idat[3]);
  assign instr_tile_rsci_d_37_33_mx0 = MUX_v_5_2_2(instr_tile_rsci_d_26_22_mx0, (tile_size_int_sva_9[4:0]),
      loops_relevancy_rsci_idat[3]);
  assign tile_size_int_lpi_1_dfm_10_5_1 = MUX_v_6_2_2(6'b000000, (tile_size_int_sva_6[10:5]),
      (loops_relevancy_rsci_idat[0]));
  assign instr_tile_rsci_d_32_27_mx0 = MUX_v_6_2_2(instr_tile_rsci_d_21_16_mx0, (tile_size_int_sva_8[10:5]),
      loops_relevancy_rsci_idat[2]);
  assign instr_tile_rsci_d_26_22_mx0 = MUX_v_5_2_2(instr_tile_rsci_d_15_11_mx0, (tile_size_int_sva_8[4:0]),
      loops_relevancy_rsci_idat[2]);
  assign instr_tile_rsci_d_21_16_mx0 = MUX_v_6_2_2(tile_size_int_lpi_1_dfm_10_5_1,
      (tile_size_int_sva_7[10:5]), loops_relevancy_rsci_idat[1]);
  assign instr_tile_rsci_d_15_11_mx0 = MUX_v_5_2_2(instr_tile_rsci_d_4_0_mx0, (tile_size_int_sva_7[4:0]),
      loops_relevancy_rsci_idat[1]);
  assign nl_tile_size_int_sva_6 = (tile_size_in_rsci_idat[4:0]) * (loops_bound_rsci_idat[10:0]);
  assign tile_size_int_sva_6 = nl_tile_size_int_sva_6[10:0];
  assign nl_tile_size_int_sva_7 = ({tile_size_int_lpi_1_dfm_10_5_1 , instr_tile_rsci_d_4_0_mx0})
      * (loops_bound_rsci_idat[21:11]);
  assign tile_size_int_sva_7 = nl_tile_size_int_sva_7[10:0];
  assign nl_tile_size_int_sva_8 = ({instr_tile_rsci_d_21_16_mx0 , instr_tile_rsci_d_15_11_mx0})
      * (loops_bound_rsci_idat[32:22]);
  assign tile_size_int_sva_8 = nl_tile_size_int_sva_8[10:0];
  assign nl_tile_size_int_sva_9 = ({instr_tile_rsci_d_32_27_mx0 , instr_tile_rsci_d_26_22_mx0})
      * (loops_bound_rsci_idat[43:33]);
  assign tile_size_int_sva_9 = nl_tile_size_int_sva_9[10:0];
  assign nl_tile_size_int_sva_10 = ({instr_tile_rsci_d_43_38_mx0 , instr_tile_rsci_d_37_33_mx0})
      * (loops_bound_rsci_idat[54:44]);
  assign tile_size_int_sva_10 = nl_tile_size_int_sva_10[10:0];
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      reg_tile_size_out_rsci_d_10_5_cse <= 6'b000000;
      reg_tile_size_out_rsci_d_4_0_cse <= 5'b00000;
      instr_tile_rsci_d_10_5 <= 6'b000000;
    end
    else if ( tile_size_and_cse ) begin
      reg_tile_size_out_rsci_d_10_5_cse <= MUX_v_6_2_2(instr_tile_rsci_d_43_38_mx0,
          (tile_size_int_sva_10[10:5]), loops_relevancy_rsci_idat[4]);
      reg_tile_size_out_rsci_d_4_0_cse <= MUX_v_5_2_2(instr_tile_rsci_d_37_33_mx0,
          (tile_size_int_sva_10[4:0]), loops_relevancy_rsci_idat[4]);
      instr_tile_rsci_d_10_5 <= tile_size_int_lpi_1_dfm_10_5_1;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      instr_bound_rsci_d_54_44 <= 11'b00000000000;
      instr_bound_rsci_d_10_0 <= 11'b00000000000;
      instr_bound_rsci_d_43_33 <= 11'b00000000000;
      instr_bound_rsci_d_21_11 <= 11'b00000000000;
      instr_bound_rsci_d_32_22 <= 11'b00000000000;
      instr_tile_rsci_d_4_0 <= 5'b00000;
      instr_tile_rsci_d_43_38 <= 6'b000000;
      instr_tile_rsci_d_37_33 <= 5'b00000;
      instr_tile_rsci_d_32_27 <= 6'b000000;
      instr_tile_rsci_d_26_22 <= 5'b00000;
      instr_tile_rsci_d_21_16 <= 6'b000000;
      instr_tile_rsci_d_15_11 <= 5'b00000;
    end
    else if ( ccs_ccore_en ) begin
      instr_bound_rsci_d_54_44 <= MUX_v_11_2_2((loops_bound_rsci_idat[54:44]), 11'b00000000001,
          loops_relevancy_rsci_idat[4]);
      instr_bound_rsci_d_10_0 <= MUX_v_11_2_2((loops_bound_rsci_idat[10:0]), 11'b00000000001,
          loops_relevancy_rsci_idat[0]);
      instr_bound_rsci_d_43_33 <= MUX_v_11_2_2((loops_bound_rsci_idat[43:33]), 11'b00000000001,
          loops_relevancy_rsci_idat[3]);
      instr_bound_rsci_d_21_11 <= MUX_v_11_2_2((loops_bound_rsci_idat[21:11]), 11'b00000000001,
          loops_relevancy_rsci_idat[1]);
      instr_bound_rsci_d_32_22 <= MUX_v_11_2_2((loops_bound_rsci_idat[32:22]), 11'b00000000001,
          loops_relevancy_rsci_idat[2]);
      instr_tile_rsci_d_4_0 <= instr_tile_rsci_d_4_0_mx0;
      instr_tile_rsci_d_43_38 <= instr_tile_rsci_d_43_38_mx0;
      instr_tile_rsci_d_37_33 <= instr_tile_rsci_d_37_33_mx0;
      instr_tile_rsci_d_32_27 <= instr_tile_rsci_d_32_27_mx0;
      instr_tile_rsci_d_26_22 <= instr_tile_rsci_d_26_22_mx0;
      instr_tile_rsci_d_21_16 <= instr_tile_rsci_d_21_16_mx0;
      instr_tile_rsci_d_15_11 <= instr_tile_rsci_d_15_11_mx0;
    end
  end

  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    tiling_unit_5_W_addr_type_L2
// ------------------------------------------------------------------


module tiling_unit_5_W_addr_type_L2 (
  loops_bound_rsc_dat, loops_relevancy_rsc_dat, tile_size_in_rsc_dat, tile_size_out_rsc_z,
      instr_bound_rsc_z, instr_tile_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [54:0] loops_bound_rsc_dat;
  input [4:0] loops_relevancy_rsc_dat;
  input [10:0] tile_size_in_rsc_dat;
  output [10:0] tile_size_out_rsc_z;
  output [54:0] instr_bound_rsc_z;
  output [54:0] instr_tile_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  tiling_unit_5_W_addr_type_L2_run tiling_unit_5_W_addr_type_L2_run_inst (
      .loops_bound_rsc_dat(loops_bound_rsc_dat),
      .loops_relevancy_rsc_dat(loops_relevancy_rsc_dat),
      .tile_size_in_rsc_dat(tile_size_in_rsc_dat),
      .tile_size_out_rsc_z(tile_size_out_rsc_z),
      .instr_bound_rsc_z(instr_bound_rsc_z),
      .instr_tile_rsc_z(instr_tile_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/tiling_unit_5_O_addr_type_L3__c8ceb417654e4d4104a4e020121ae510b7ce_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   r0678912@amazone.esat.kuleuven.be
//  Generated date: Tue Jul 13 10:57:58 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    tiling_unit_5_O_addr_type_L3_run
// ------------------------------------------------------------------


module tiling_unit_5_O_addr_type_L3_run (
  loops_bound_rsc_dat, loops_relevancy_rsc_dat, tile_size_in_rsc_dat, tile_size_out_rsc_z,
      instr_bound_rsc_z, instr_tile_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [69:0] loops_bound_rsc_dat;
  input [4:0] loops_relevancy_rsc_dat;
  input [13:0] tile_size_in_rsc_dat;
  output [13:0] tile_size_out_rsc_z;
  output [69:0] instr_bound_rsc_z;
  output [69:0] instr_tile_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [69:0] loops_bound_rsci_idat;
  wire [4:0] loops_relevancy_rsci_idat;
  wire [13:0] tile_size_in_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [13:0] instr_bound_rsci_d_69_56;
  reg [13:0] instr_bound_rsci_d_55_42;
  reg [13:0] instr_bound_rsci_d_41_28;
  reg [13:0] instr_bound_rsci_d_27_14;
  reg [13:0] instr_bound_rsci_d_13_0;
  reg [4:0] instr_tile_rsci_d_13_9;
  reg [8:0] instr_tile_rsci_d_8_0;
  reg [4:0] instr_tile_rsci_d_55_51;
  reg [8:0] instr_tile_rsci_d_50_42;
  reg [4:0] instr_tile_rsci_d_41_37;
  reg [8:0] instr_tile_rsci_d_36_28;
  reg [4:0] instr_tile_rsci_d_27_23;
  reg [8:0] instr_tile_rsci_d_22_14;
  reg [4:0] reg_tile_size_out_rsci_d_13_9_cse;
  reg [8:0] reg_tile_size_out_rsci_d_8_0_cse;
  wire [8:0] instr_tile_rsci_d_8_0_mx0;
  wire [4:0] instr_tile_rsci_d_55_51_mx0;
  wire [8:0] instr_tile_rsci_d_50_42_mx0;
  wire [4:0] tile_size_int_lpi_1_dfm_13_9_1;
  wire [4:0] instr_tile_rsci_d_41_37_mx0;
  wire [8:0] instr_tile_rsci_d_36_28_mx0;
  wire [4:0] instr_tile_rsci_d_27_23_mx0;
  wire [8:0] instr_tile_rsci_d_22_14_mx0;
  wire [13:0] tile_size_int_sva_6;
  wire [22:0] nl_tile_size_int_sva_6;
  wire [13:0] tile_size_int_sva_7;
  wire [27:0] nl_tile_size_int_sva_7;
  wire [13:0] tile_size_int_sva_8;
  wire [27:0] nl_tile_size_int_sva_8;
  wire [13:0] tile_size_int_sva_9;
  wire [27:0] nl_tile_size_int_sva_9;
  wire [13:0] tile_size_int_sva_10;
  wire [27:0] nl_tile_size_int_sva_10;
  wire tile_size_and_cse;


  // Interconnect Declarations for Component Instantiations 
  wire [69:0] nl_instr_bound_rsci_d;
  assign nl_instr_bound_rsci_d = {instr_bound_rsci_d_69_56 , instr_bound_rsci_d_55_42
      , instr_bound_rsci_d_41_28 , instr_bound_rsci_d_27_14 , instr_bound_rsci_d_13_0};
  wire [69:0] nl_instr_tile_rsci_d;
  assign nl_instr_tile_rsci_d = {reg_tile_size_out_rsci_d_13_9_cse , reg_tile_size_out_rsci_d_8_0_cse
      , instr_tile_rsci_d_55_51 , instr_tile_rsci_d_50_42 , instr_tile_rsci_d_41_37
      , instr_tile_rsci_d_36_28 , instr_tile_rsci_d_27_23 , instr_tile_rsci_d_22_14
      , instr_tile_rsci_d_13_9 , instr_tile_rsci_d_8_0};
  wire [13:0] nl_tile_size_out_rsci_d;
  assign nl_tile_size_out_rsci_d = {reg_tile_size_out_rsci_d_13_9_cse , reg_tile_size_out_rsci_d_8_0_cse};
  ccs_in_v1 #(.rscid(32'sd11),
  .width(32'sd70)) loops_bound_rsci (
      .dat(loops_bound_rsc_dat),
      .idat(loops_bound_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd12),
  .width(32'sd5)) loops_relevancy_rsci (
      .dat(loops_relevancy_rsc_dat),
      .idat(loops_relevancy_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd14),
  .width(32'sd70)) instr_bound_rsci (
      .d(nl_instr_bound_rsci_d[69:0]),
      .z(instr_bound_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd15),
  .width(32'sd70)) instr_tile_rsci (
      .d(nl_instr_tile_rsci_d[69:0]),
      .z(instr_tile_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd126),
  .width(32'sd14)) tile_size_in_rsci (
      .dat(tile_size_in_rsc_dat),
      .idat(tile_size_in_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd127),
  .width(32'sd14)) tile_size_out_rsci (
      .d(nl_tile_size_out_rsci_d[13:0]),
      .z(tile_size_out_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd135),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign tile_size_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  assign instr_tile_rsci_d_8_0_mx0 = MUX_v_9_2_2((tile_size_in_rsci_idat[8:0]), (tile_size_int_sva_6[8:0]),
      loops_relevancy_rsci_idat[0]);
  assign instr_tile_rsci_d_55_51_mx0 = MUX_v_5_2_2(instr_tile_rsci_d_41_37_mx0, (tile_size_int_sva_9[13:9]),
      loops_relevancy_rsci_idat[3]);
  assign instr_tile_rsci_d_50_42_mx0 = MUX_v_9_2_2(instr_tile_rsci_d_36_28_mx0, (tile_size_int_sva_9[8:0]),
      loops_relevancy_rsci_idat[3]);
  assign tile_size_int_lpi_1_dfm_13_9_1 = MUX_v_5_2_2(5'b00000, (tile_size_int_sva_6[13:9]),
      (loops_relevancy_rsci_idat[0]));
  assign instr_tile_rsci_d_41_37_mx0 = MUX_v_5_2_2(instr_tile_rsci_d_27_23_mx0, (tile_size_int_sva_8[13:9]),
      loops_relevancy_rsci_idat[2]);
  assign instr_tile_rsci_d_36_28_mx0 = MUX_v_9_2_2(instr_tile_rsci_d_22_14_mx0, (tile_size_int_sva_8[8:0]),
      loops_relevancy_rsci_idat[2]);
  assign instr_tile_rsci_d_27_23_mx0 = MUX_v_5_2_2(tile_size_int_lpi_1_dfm_13_9_1,
      (tile_size_int_sva_7[13:9]), loops_relevancy_rsci_idat[1]);
  assign instr_tile_rsci_d_22_14_mx0 = MUX_v_9_2_2(instr_tile_rsci_d_8_0_mx0, (tile_size_int_sva_7[8:0]),
      loops_relevancy_rsci_idat[1]);
  assign nl_tile_size_int_sva_6 = (tile_size_in_rsci_idat[8:0]) * (loops_bound_rsci_idat[13:0]);
  assign tile_size_int_sva_6 = nl_tile_size_int_sva_6[13:0];
  assign nl_tile_size_int_sva_7 = ({tile_size_int_lpi_1_dfm_13_9_1 , instr_tile_rsci_d_8_0_mx0})
      * (loops_bound_rsci_idat[27:14]);
  assign tile_size_int_sva_7 = nl_tile_size_int_sva_7[13:0];
  assign nl_tile_size_int_sva_8 = ({instr_tile_rsci_d_27_23_mx0 , instr_tile_rsci_d_22_14_mx0})
      * (loops_bound_rsci_idat[41:28]);
  assign tile_size_int_sva_8 = nl_tile_size_int_sva_8[13:0];
  assign nl_tile_size_int_sva_9 = ({instr_tile_rsci_d_41_37_mx0 , instr_tile_rsci_d_36_28_mx0})
      * (loops_bound_rsci_idat[55:42]);
  assign tile_size_int_sva_9 = nl_tile_size_int_sva_9[13:0];
  assign nl_tile_size_int_sva_10 = ({instr_tile_rsci_d_55_51_mx0 , instr_tile_rsci_d_50_42_mx0})
      * (loops_bound_rsci_idat[69:56]);
  assign tile_size_int_sva_10 = nl_tile_size_int_sva_10[13:0];
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      reg_tile_size_out_rsci_d_13_9_cse <= 5'b00000;
      reg_tile_size_out_rsci_d_8_0_cse <= 9'b000000000;
      instr_tile_rsci_d_13_9 <= 5'b00000;
    end
    else if ( tile_size_and_cse ) begin
      reg_tile_size_out_rsci_d_13_9_cse <= MUX_v_5_2_2(instr_tile_rsci_d_55_51_mx0,
          (tile_size_int_sva_10[13:9]), loops_relevancy_rsci_idat[4]);
      reg_tile_size_out_rsci_d_8_0_cse <= MUX_v_9_2_2(instr_tile_rsci_d_50_42_mx0,
          (tile_size_int_sva_10[8:0]), loops_relevancy_rsci_idat[4]);
      instr_tile_rsci_d_13_9 <= tile_size_int_lpi_1_dfm_13_9_1;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      instr_bound_rsci_d_69_56 <= 14'b00000000000000;
      instr_bound_rsci_d_13_0 <= 14'b00000000000000;
      instr_bound_rsci_d_55_42 <= 14'b00000000000000;
      instr_bound_rsci_d_27_14 <= 14'b00000000000000;
      instr_bound_rsci_d_41_28 <= 14'b00000000000000;
      instr_tile_rsci_d_8_0 <= 9'b000000000;
      instr_tile_rsci_d_55_51 <= 5'b00000;
      instr_tile_rsci_d_50_42 <= 9'b000000000;
      instr_tile_rsci_d_41_37 <= 5'b00000;
      instr_tile_rsci_d_36_28 <= 9'b000000000;
      instr_tile_rsci_d_27_23 <= 5'b00000;
      instr_tile_rsci_d_22_14 <= 9'b000000000;
    end
    else if ( ccs_ccore_en ) begin
      instr_bound_rsci_d_69_56 <= MUX_v_14_2_2((loops_bound_rsci_idat[69:56]), 14'b00000000000001,
          loops_relevancy_rsci_idat[4]);
      instr_bound_rsci_d_13_0 <= MUX_v_14_2_2((loops_bound_rsci_idat[13:0]), 14'b00000000000001,
          loops_relevancy_rsci_idat[0]);
      instr_bound_rsci_d_55_42 <= MUX_v_14_2_2((loops_bound_rsci_idat[55:42]), 14'b00000000000001,
          loops_relevancy_rsci_idat[3]);
      instr_bound_rsci_d_27_14 <= MUX_v_14_2_2((loops_bound_rsci_idat[27:14]), 14'b00000000000001,
          loops_relevancy_rsci_idat[1]);
      instr_bound_rsci_d_41_28 <= MUX_v_14_2_2((loops_bound_rsci_idat[41:28]), 14'b00000000000001,
          loops_relevancy_rsci_idat[2]);
      instr_tile_rsci_d_8_0 <= instr_tile_rsci_d_8_0_mx0;
      instr_tile_rsci_d_55_51 <= instr_tile_rsci_d_55_51_mx0;
      instr_tile_rsci_d_50_42 <= instr_tile_rsci_d_50_42_mx0;
      instr_tile_rsci_d_41_37 <= instr_tile_rsci_d_41_37_mx0;
      instr_tile_rsci_d_36_28 <= instr_tile_rsci_d_36_28_mx0;
      instr_tile_rsci_d_27_23 <= instr_tile_rsci_d_27_23_mx0;
      instr_tile_rsci_d_22_14 <= instr_tile_rsci_d_22_14_mx0;
    end
  end

  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [0:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    tiling_unit_5_O_addr_type_L3
// ------------------------------------------------------------------


module tiling_unit_5_O_addr_type_L3 (
  loops_bound_rsc_dat, loops_relevancy_rsc_dat, tile_size_in_rsc_dat, tile_size_out_rsc_z,
      instr_bound_rsc_z, instr_tile_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [69:0] loops_bound_rsc_dat;
  input [4:0] loops_relevancy_rsc_dat;
  input [13:0] tile_size_in_rsc_dat;
  output [13:0] tile_size_out_rsc_z;
  output [69:0] instr_bound_rsc_z;
  output [69:0] instr_tile_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  tiling_unit_5_O_addr_type_L3_run tiling_unit_5_O_addr_type_L3_run_inst (
      .loops_bound_rsc_dat(loops_bound_rsc_dat),
      .loops_relevancy_rsc_dat(loops_relevancy_rsc_dat),
      .tile_size_in_rsc_dat(tile_size_in_rsc_dat),
      .tile_size_out_rsc_z(tile_size_out_rsc_z),
      .instr_bound_rsc_z(instr_bound_rsc_z),
      .instr_tile_rsc_z(instr_tile_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/tiling_unit_5_O_addr_type_L2__62fbec45f0c0ed28ff5c917a6fb9ea42b629_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   r0678912@amazone.esat.kuleuven.be
//  Generated date: Tue Jul 13 10:58:00 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    tiling_unit_5_O_addr_type_L2_run
// ------------------------------------------------------------------


module tiling_unit_5_O_addr_type_L2_run (
  loops_bound_rsc_dat, loops_relevancy_rsc_dat, tile_size_in_rsc_dat, tile_size_out_rsc_z,
      instr_bound_rsc_z, instr_tile_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [44:0] loops_bound_rsc_dat;
  input [4:0] loops_relevancy_rsc_dat;
  input [8:0] tile_size_in_rsc_dat;
  output [8:0] tile_size_out_rsc_z;
  output [44:0] instr_bound_rsc_z;
  output [44:0] instr_tile_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [44:0] loops_bound_rsci_idat;
  wire [4:0] loops_relevancy_rsci_idat;
  wire [8:0] tile_size_in_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [8:0] instr_bound_rsci_d_44_36;
  reg [8:0] instr_bound_rsci_d_35_27;
  reg [8:0] instr_bound_rsci_d_26_18;
  reg [8:0] instr_bound_rsci_d_17_9;
  reg [8:0] instr_bound_rsci_d_8_0;
  reg [3:0] instr_tile_rsci_d_8_5;
  reg [4:0] instr_tile_rsci_d_4_0;
  reg [3:0] instr_tile_rsci_d_35_32;
  reg [4:0] instr_tile_rsci_d_31_27;
  reg [3:0] instr_tile_rsci_d_26_23;
  reg [4:0] instr_tile_rsci_d_22_18;
  reg [3:0] instr_tile_rsci_d_17_14;
  reg [4:0] instr_tile_rsci_d_13_9;
  reg [3:0] reg_tile_size_out_rsci_d_8_5_cse;
  reg [4:0] reg_tile_size_out_rsci_d_4_0_cse;
  wire [4:0] instr_tile_rsci_d_4_0_mx0;
  wire [3:0] instr_tile_rsci_d_35_32_mx0;
  wire [4:0] instr_tile_rsci_d_31_27_mx0;
  wire [3:0] tile_size_int_lpi_1_dfm_8_5_1;
  wire [3:0] instr_tile_rsci_d_26_23_mx0;
  wire [4:0] instr_tile_rsci_d_22_18_mx0;
  wire [3:0] instr_tile_rsci_d_17_14_mx0;
  wire [4:0] instr_tile_rsci_d_13_9_mx0;
  wire [8:0] tile_size_int_sva_6;
  wire [13:0] nl_tile_size_int_sva_6;
  wire [8:0] tile_size_int_sva_7;
  wire [17:0] nl_tile_size_int_sva_7;
  wire [8:0] tile_size_int_sva_8;
  wire [17:0] nl_tile_size_int_sva_8;
  wire [8:0] tile_size_int_sva_9;
  wire [17:0] nl_tile_size_int_sva_9;
  wire [8:0] tile_size_int_sva_10;
  wire [17:0] nl_tile_size_int_sva_10;
  wire tile_size_and_cse;


  // Interconnect Declarations for Component Instantiations 
  wire [44:0] nl_instr_bound_rsci_d;
  assign nl_instr_bound_rsci_d = {instr_bound_rsci_d_44_36 , instr_bound_rsci_d_35_27
      , instr_bound_rsci_d_26_18 , instr_bound_rsci_d_17_9 , instr_bound_rsci_d_8_0};
  wire [44:0] nl_instr_tile_rsci_d;
  assign nl_instr_tile_rsci_d = {reg_tile_size_out_rsci_d_8_5_cse , reg_tile_size_out_rsci_d_4_0_cse
      , instr_tile_rsci_d_35_32 , instr_tile_rsci_d_31_27 , instr_tile_rsci_d_26_23
      , instr_tile_rsci_d_22_18 , instr_tile_rsci_d_17_14 , instr_tile_rsci_d_13_9
      , instr_tile_rsci_d_8_5 , instr_tile_rsci_d_4_0};
  wire [8:0] nl_tile_size_out_rsci_d;
  assign nl_tile_size_out_rsci_d = {reg_tile_size_out_rsci_d_8_5_cse , reg_tile_size_out_rsci_d_4_0_cse};
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd45)) loops_bound_rsci (
      .dat(loops_bound_rsc_dat),
      .idat(loops_bound_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd7),
  .width(32'sd5)) loops_relevancy_rsci (
      .dat(loops_relevancy_rsc_dat),
      .idat(loops_relevancy_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd9),
  .width(32'sd45)) instr_bound_rsci (
      .d(nl_instr_bound_rsci_d[44:0]),
      .z(instr_bound_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd10),
  .width(32'sd45)) instr_tile_rsci (
      .d(nl_instr_tile_rsci_d[44:0]),
      .z(instr_tile_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd128),
  .width(32'sd9)) tile_size_in_rsci (
      .dat(tile_size_in_rsc_dat),
      .idat(tile_size_in_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd129),
  .width(32'sd9)) tile_size_out_rsci (
      .d(nl_tile_size_out_rsci_d[8:0]),
      .z(tile_size_out_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd136),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign tile_size_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  assign instr_tile_rsci_d_4_0_mx0 = MUX_v_5_2_2((tile_size_in_rsci_idat[4:0]), (tile_size_int_sva_6[4:0]),
      loops_relevancy_rsci_idat[0]);
  assign instr_tile_rsci_d_35_32_mx0 = MUX_v_4_2_2(instr_tile_rsci_d_26_23_mx0, (tile_size_int_sva_9[8:5]),
      loops_relevancy_rsci_idat[3]);
  assign instr_tile_rsci_d_31_27_mx0 = MUX_v_5_2_2(instr_tile_rsci_d_22_18_mx0, (tile_size_int_sva_9[4:0]),
      loops_relevancy_rsci_idat[3]);
  assign tile_size_int_lpi_1_dfm_8_5_1 = MUX_v_4_2_2(4'b0000, (tile_size_int_sva_6[8:5]),
      (loops_relevancy_rsci_idat[0]));
  assign instr_tile_rsci_d_26_23_mx0 = MUX_v_4_2_2(instr_tile_rsci_d_17_14_mx0, (tile_size_int_sva_8[8:5]),
      loops_relevancy_rsci_idat[2]);
  assign instr_tile_rsci_d_22_18_mx0 = MUX_v_5_2_2(instr_tile_rsci_d_13_9_mx0, (tile_size_int_sva_8[4:0]),
      loops_relevancy_rsci_idat[2]);
  assign instr_tile_rsci_d_17_14_mx0 = MUX_v_4_2_2(tile_size_int_lpi_1_dfm_8_5_1,
      (tile_size_int_sva_7[8:5]), loops_relevancy_rsci_idat[1]);
  assign instr_tile_rsci_d_13_9_mx0 = MUX_v_5_2_2(instr_tile_rsci_d_4_0_mx0, (tile_size_int_sva_7[4:0]),
      loops_relevancy_rsci_idat[1]);
  assign nl_tile_size_int_sva_6 = (tile_size_in_rsci_idat[4:0]) * (loops_bound_rsci_idat[8:0]);
  assign tile_size_int_sva_6 = nl_tile_size_int_sva_6[8:0];
  assign nl_tile_size_int_sva_7 = ({tile_size_int_lpi_1_dfm_8_5_1 , instr_tile_rsci_d_4_0_mx0})
      * (loops_bound_rsci_idat[17:9]);
  assign tile_size_int_sva_7 = nl_tile_size_int_sva_7[8:0];
  assign nl_tile_size_int_sva_8 = ({instr_tile_rsci_d_17_14_mx0 , instr_tile_rsci_d_13_9_mx0})
      * (loops_bound_rsci_idat[26:18]);
  assign tile_size_int_sva_8 = nl_tile_size_int_sva_8[8:0];
  assign nl_tile_size_int_sva_9 = ({instr_tile_rsci_d_26_23_mx0 , instr_tile_rsci_d_22_18_mx0})
      * (loops_bound_rsci_idat[35:27]);
  assign tile_size_int_sva_9 = nl_tile_size_int_sva_9[8:0];
  assign nl_tile_size_int_sva_10 = ({instr_tile_rsci_d_35_32_mx0 , instr_tile_rsci_d_31_27_mx0})
      * (loops_bound_rsci_idat[44:36]);
  assign tile_size_int_sva_10 = nl_tile_size_int_sva_10[8:0];
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      reg_tile_size_out_rsci_d_8_5_cse <= 4'b0000;
      reg_tile_size_out_rsci_d_4_0_cse <= 5'b00000;
      instr_tile_rsci_d_8_5 <= 4'b0000;
    end
    else if ( tile_size_and_cse ) begin
      reg_tile_size_out_rsci_d_8_5_cse <= MUX_v_4_2_2(instr_tile_rsci_d_35_32_mx0,
          (tile_size_int_sva_10[8:5]), loops_relevancy_rsci_idat[4]);
      reg_tile_size_out_rsci_d_4_0_cse <= MUX_v_5_2_2(instr_tile_rsci_d_31_27_mx0,
          (tile_size_int_sva_10[4:0]), loops_relevancy_rsci_idat[4]);
      instr_tile_rsci_d_8_5 <= tile_size_int_lpi_1_dfm_8_5_1;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      instr_bound_rsci_d_44_36 <= 9'b000000000;
      instr_bound_rsci_d_8_0 <= 9'b000000000;
      instr_bound_rsci_d_35_27 <= 9'b000000000;
      instr_bound_rsci_d_17_9 <= 9'b000000000;
      instr_bound_rsci_d_26_18 <= 9'b000000000;
      instr_tile_rsci_d_4_0 <= 5'b00000;
      instr_tile_rsci_d_35_32 <= 4'b0000;
      instr_tile_rsci_d_31_27 <= 5'b00000;
      instr_tile_rsci_d_26_23 <= 4'b0000;
      instr_tile_rsci_d_22_18 <= 5'b00000;
      instr_tile_rsci_d_17_14 <= 4'b0000;
      instr_tile_rsci_d_13_9 <= 5'b00000;
    end
    else if ( ccs_ccore_en ) begin
      instr_bound_rsci_d_44_36 <= MUX_v_9_2_2((loops_bound_rsci_idat[44:36]), 9'b000000001,
          loops_relevancy_rsci_idat[4]);
      instr_bound_rsci_d_8_0 <= MUX_v_9_2_2((loops_bound_rsci_idat[8:0]), 9'b000000001,
          loops_relevancy_rsci_idat[0]);
      instr_bound_rsci_d_35_27 <= MUX_v_9_2_2((loops_bound_rsci_idat[35:27]), 9'b000000001,
          loops_relevancy_rsci_idat[3]);
      instr_bound_rsci_d_17_9 <= MUX_v_9_2_2((loops_bound_rsci_idat[17:9]), 9'b000000001,
          loops_relevancy_rsci_idat[1]);
      instr_bound_rsci_d_26_18 <= MUX_v_9_2_2((loops_bound_rsci_idat[26:18]), 9'b000000001,
          loops_relevancy_rsci_idat[2]);
      instr_tile_rsci_d_4_0 <= instr_tile_rsci_d_4_0_mx0;
      instr_tile_rsci_d_35_32 <= instr_tile_rsci_d_35_32_mx0;
      instr_tile_rsci_d_31_27 <= instr_tile_rsci_d_31_27_mx0;
      instr_tile_rsci_d_26_23 <= instr_tile_rsci_d_26_23_mx0;
      instr_tile_rsci_d_22_18 <= instr_tile_rsci_d_22_18_mx0;
      instr_tile_rsci_d_17_14 <= instr_tile_rsci_d_17_14_mx0;
      instr_tile_rsci_d_13_9 <= instr_tile_rsci_d_13_9_mx0;
    end
  end

  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    tiling_unit_5_O_addr_type_L2
// ------------------------------------------------------------------


module tiling_unit_5_O_addr_type_L2 (
  loops_bound_rsc_dat, loops_relevancy_rsc_dat, tile_size_in_rsc_dat, tile_size_out_rsc_z,
      instr_bound_rsc_z, instr_tile_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [44:0] loops_bound_rsc_dat;
  input [4:0] loops_relevancy_rsc_dat;
  input [8:0] tile_size_in_rsc_dat;
  output [8:0] tile_size_out_rsc_z;
  output [44:0] instr_bound_rsc_z;
  output [44:0] instr_tile_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  tiling_unit_5_O_addr_type_L2_run tiling_unit_5_O_addr_type_L2_run_inst (
      .loops_bound_rsc_dat(loops_bound_rsc_dat),
      .loops_relevancy_rsc_dat(loops_relevancy_rsc_dat),
      .tile_size_in_rsc_dat(tile_size_in_rsc_dat),
      .tile_size_out_rsc_z(tile_size_out_rsc_z),
      .instr_bound_rsc_z(instr_bound_rsc_z),
      .instr_tile_rsc_z(instr_tile_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/tiling_unit_5_O_addr_type_L1__8602e08520fb27a65174dadf7fa1b550aec7_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   r0678912@amazone.esat.kuleuven.be
//  Generated date: Tue Jul 13 10:58:02 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    tiling_unit_5_O_addr_type_L1_run
// ------------------------------------------------------------------


module tiling_unit_5_O_addr_type_L1_run (
  loops_bound_rsc_dat, loops_relevancy_rsc_dat, tile_size_in_rsc_dat, tile_size_out_rsc_z,
      instr_bound_rsc_z, instr_tile_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [24:0] loops_bound_rsc_dat;
  input [4:0] loops_relevancy_rsc_dat;
  input [4:0] tile_size_in_rsc_dat;
  output [4:0] tile_size_out_rsc_z;
  output [24:0] instr_bound_rsc_z;
  output [24:0] instr_tile_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [24:0] loops_bound_rsci_idat;
  wire [4:0] loops_relevancy_rsci_idat;
  wire [4:0] tile_size_in_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [4:0] instr_bound_rsci_d_24_20;
  reg [4:0] instr_bound_rsci_d_19_15;
  reg [4:0] instr_bound_rsci_d_14_10;
  reg [4:0] instr_bound_rsci_d_9_5;
  reg [4:0] instr_bound_rsci_d_4_0;
  reg [4:0] instr_tile_rsci_d_19_15;
  reg [4:0] instr_tile_rsci_d_14_10;
  reg [4:0] instr_tile_rsci_d_9_5;
  reg [4:0] instr_tile_rsci_d_4_0;
  reg [4:0] reg_tile_size_out_rsci_d_cse;
  wire [4:0] instr_tile_rsci_d_4_0_mx0;
  wire [4:0] instr_tile_rsci_d_19_15_mx0;
  wire [4:0] instr_tile_rsci_d_9_5_mx0;
  wire [4:0] instr_tile_rsci_d_14_10_mx0;
  wire tile_size_and_cse;

  wire[4:0] for_5_if_mul_nl;
  wire[9:0] nl_for_5_if_mul_nl;
  wire[4:0] for_1_if_mul_nl;
  wire[9:0] nl_for_1_if_mul_nl;
  wire[4:0] for_4_if_mul_nl;
  wire[9:0] nl_for_4_if_mul_nl;
  wire[4:0] for_2_if_mul_nl;
  wire[9:0] nl_for_2_if_mul_nl;
  wire[4:0] for_3_if_mul_nl;
  wire[9:0] nl_for_3_if_mul_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [24:0] nl_instr_bound_rsci_d;
  assign nl_instr_bound_rsci_d = {instr_bound_rsci_d_24_20 , instr_bound_rsci_d_19_15
      , instr_bound_rsci_d_14_10 , instr_bound_rsci_d_9_5 , instr_bound_rsci_d_4_0};
  wire [24:0] nl_instr_tile_rsci_d;
  assign nl_instr_tile_rsci_d = {reg_tile_size_out_rsci_d_cse , instr_tile_rsci_d_19_15
      , instr_tile_rsci_d_14_10 , instr_tile_rsci_d_9_5 , instr_tile_rsci_d_4_0};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd25)) loops_bound_rsci (
      .dat(loops_bound_rsc_dat),
      .idat(loops_bound_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd5)) loops_relevancy_rsci (
      .dat(loops_relevancy_rsc_dat),
      .idat(loops_relevancy_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd4),
  .width(32'sd25)) instr_bound_rsci (
      .d(nl_instr_bound_rsci_d[24:0]),
      .z(instr_bound_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd5),
  .width(32'sd25)) instr_tile_rsci (
      .d(nl_instr_tile_rsci_d[24:0]),
      .z(instr_tile_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd130),
  .width(32'sd5)) tile_size_in_rsci (
      .dat(tile_size_in_rsc_dat),
      .idat(tile_size_in_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd131),
  .width(32'sd5)) tile_size_out_rsci (
      .d(reg_tile_size_out_rsci_d_cse),
      .z(tile_size_out_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd137),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign tile_size_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  assign nl_for_1_if_mul_nl = tile_size_in_rsci_idat * (loops_bound_rsci_idat[4:0]);
  assign for_1_if_mul_nl = nl_for_1_if_mul_nl[4:0];
  assign instr_tile_rsci_d_4_0_mx0 = MUX_v_5_2_2(tile_size_in_rsci_idat, for_1_if_mul_nl,
      loops_relevancy_rsci_idat[0]);
  assign nl_for_4_if_mul_nl = instr_tile_rsci_d_14_10_mx0 * (loops_bound_rsci_idat[19:15]);
  assign for_4_if_mul_nl = nl_for_4_if_mul_nl[4:0];
  assign instr_tile_rsci_d_19_15_mx0 = MUX_v_5_2_2(instr_tile_rsci_d_14_10_mx0, for_4_if_mul_nl,
      loops_relevancy_rsci_idat[3]);
  assign nl_for_2_if_mul_nl = instr_tile_rsci_d_4_0_mx0 * (loops_bound_rsci_idat[9:5]);
  assign for_2_if_mul_nl = nl_for_2_if_mul_nl[4:0];
  assign instr_tile_rsci_d_9_5_mx0 = MUX_v_5_2_2(instr_tile_rsci_d_4_0_mx0, for_2_if_mul_nl,
      loops_relevancy_rsci_idat[1]);
  assign nl_for_3_if_mul_nl = instr_tile_rsci_d_9_5_mx0 * (loops_bound_rsci_idat[14:10]);
  assign for_3_if_mul_nl = nl_for_3_if_mul_nl[4:0];
  assign instr_tile_rsci_d_14_10_mx0 = MUX_v_5_2_2(instr_tile_rsci_d_9_5_mx0, for_3_if_mul_nl,
      loops_relevancy_rsci_idat[2]);
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      reg_tile_size_out_rsci_d_cse <= 5'b00000;
      instr_tile_rsci_d_4_0 <= 5'b00000;
      instr_tile_rsci_d_19_15 <= 5'b00000;
      instr_tile_rsci_d_9_5 <= 5'b00000;
      instr_tile_rsci_d_14_10 <= 5'b00000;
    end
    else if ( tile_size_and_cse ) begin
      reg_tile_size_out_rsci_d_cse <= MUX_v_5_2_2(instr_tile_rsci_d_19_15_mx0, for_5_if_mul_nl,
          loops_relevancy_rsci_idat[4]);
      instr_tile_rsci_d_4_0 <= instr_tile_rsci_d_4_0_mx0;
      instr_tile_rsci_d_19_15 <= instr_tile_rsci_d_19_15_mx0;
      instr_tile_rsci_d_9_5 <= instr_tile_rsci_d_9_5_mx0;
      instr_tile_rsci_d_14_10 <= instr_tile_rsci_d_14_10_mx0;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      instr_bound_rsci_d_24_20 <= 5'b00000;
      instr_bound_rsci_d_4_0 <= 5'b00000;
      instr_bound_rsci_d_19_15 <= 5'b00000;
      instr_bound_rsci_d_9_5 <= 5'b00000;
      instr_bound_rsci_d_14_10 <= 5'b00000;
    end
    else if ( ccs_ccore_en ) begin
      instr_bound_rsci_d_24_20 <= MUX_v_5_2_2((loops_bound_rsci_idat[24:20]), 5'b00001,
          loops_relevancy_rsci_idat[4]);
      instr_bound_rsci_d_4_0 <= MUX_v_5_2_2((loops_bound_rsci_idat[4:0]), 5'b00001,
          loops_relevancy_rsci_idat[0]);
      instr_bound_rsci_d_19_15 <= MUX_v_5_2_2((loops_bound_rsci_idat[19:15]), 5'b00001,
          loops_relevancy_rsci_idat[3]);
      instr_bound_rsci_d_9_5 <= MUX_v_5_2_2((loops_bound_rsci_idat[9:5]), 5'b00001,
          loops_relevancy_rsci_idat[1]);
      instr_bound_rsci_d_14_10 <= MUX_v_5_2_2((loops_bound_rsci_idat[14:10]), 5'b00001,
          loops_relevancy_rsci_idat[2]);
    end
  end
  assign nl_for_5_if_mul_nl = instr_tile_rsci_d_19_15_mx0 * (loops_bound_rsci_idat[24:20]);
  assign for_5_if_mul_nl = nl_for_5_if_mul_nl[4:0];

  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    tiling_unit_5_O_addr_type_L1
// ------------------------------------------------------------------


module tiling_unit_5_O_addr_type_L1 (
  loops_bound_rsc_dat, loops_relevancy_rsc_dat, tile_size_in_rsc_dat, tile_size_out_rsc_z,
      instr_bound_rsc_z, instr_tile_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [24:0] loops_bound_rsc_dat;
  input [4:0] loops_relevancy_rsc_dat;
  input [4:0] tile_size_in_rsc_dat;
  output [4:0] tile_size_out_rsc_z;
  output [24:0] instr_bound_rsc_z;
  output [24:0] instr_tile_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  tiling_unit_5_O_addr_type_L1_run tiling_unit_5_O_addr_type_L1_run_inst (
      .loops_bound_rsc_dat(loops_bound_rsc_dat),
      .loops_relevancy_rsc_dat(loops_relevancy_rsc_dat),
      .tile_size_in_rsc_dat(tile_size_in_rsc_dat),
      .tile_size_out_rsc_z(tile_size_out_rsc_z),
      .instr_bound_rsc_z(instr_bound_rsc_z),
      .instr_tile_rsc_z(instr_tile_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   r0678912@amazone.esat.kuleuven.be
//  Generated date: Tue Jul 13 11:42:27 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_run_fsm
    (
  clk, rst, run_wen, fsm_output
);
  input clk;
  input rst;
  input run_wen;
  output [7:0] fsm_output;
  reg [7:0] fsm_output;


  // FSM State Type Declaration for config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_run_fsm_1
  parameter
    run_rlp_C_0 = 3'd0,
    main_C_0 = 3'd1,
    main_C_1 = 3'd2,
    main_C_2 = 3'd3,
    main_C_3 = 3'd4,
    main_C_4 = 3'd5,
    main_C_5 = 3'd6,
    main_C_6 = 3'd7;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 8'b00000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 8'b00000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 8'b00001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 8'b00010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 8'b00100000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 8'b01000000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 8'b10000000;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 8'b00000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_staller
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_staller
    (
  run_wen, layer_instruction_in_rsci_wen_comp, O_instr_L1_out_rsci_wen_comp, O_instr_L2_out_rsci_wen_comp,
      O_instr_L3_out_rsci_wen_comp, I_instr_L1_out_rsci_wen_comp, I_instr_L2_out_rsci_wen_comp,
      I_instr_L3_out_rsci_wen_comp, W_instr_L1_out_rsci_wen_comp, W_instr_L2_out_rsci_wen_comp,
      W_instr_L3_out_rsci_wen_comp
);
  output run_wen;
  input layer_instruction_in_rsci_wen_comp;
  input O_instr_L1_out_rsci_wen_comp;
  input O_instr_L2_out_rsci_wen_comp;
  input O_instr_L3_out_rsci_wen_comp;
  input I_instr_L1_out_rsci_wen_comp;
  input I_instr_L2_out_rsci_wen_comp;
  input I_instr_L3_out_rsci_wen_comp;
  input W_instr_L1_out_rsci_wen_comp;
  input W_instr_L2_out_rsci_wen_comp;
  input W_instr_L3_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = layer_instruction_in_rsci_wen_comp & O_instr_L1_out_rsci_wen_comp
      & O_instr_L2_out_rsci_wen_comp & O_instr_L3_out_rsci_wen_comp & I_instr_L1_out_rsci_wen_comp
      & I_instr_L2_out_rsci_wen_comp & I_instr_L3_out_rsci_wen_comp & W_instr_L1_out_rsci_wen_comp
      & W_instr_L2_out_rsci_wen_comp & W_instr_L3_out_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_wait_dp
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_wait_dp
    (
  ensig_cgo_iro, W_tiling_unit_L3_run_cmp_ccs_ccore_en, ensig_cgo_iro_1, W_tiling_unit_L2_run_cmp_ccs_ccore_en,
      ensig_cgo_iro_2, O_tiling_unit_L3_run_cmp_ccs_ccore_en, ensig_cgo_iro_3, O_tiling_unit_L2_run_cmp_ccs_ccore_en,
      ensig_cgo_iro_4, O_tiling_unit_L1_run_cmp_ccs_ccore_en, run_wen, ensig_cgo,
      ensig_cgo_1, ensig_cgo_2, ensig_cgo_3, ensig_cgo_4
);
  input ensig_cgo_iro;
  output W_tiling_unit_L3_run_cmp_ccs_ccore_en;
  input ensig_cgo_iro_1;
  output W_tiling_unit_L2_run_cmp_ccs_ccore_en;
  input ensig_cgo_iro_2;
  output O_tiling_unit_L3_run_cmp_ccs_ccore_en;
  input ensig_cgo_iro_3;
  output O_tiling_unit_L2_run_cmp_ccs_ccore_en;
  input ensig_cgo_iro_4;
  output O_tiling_unit_L1_run_cmp_ccs_ccore_en;
  input run_wen;
  input ensig_cgo;
  input ensig_cgo_1;
  input ensig_cgo_2;
  input ensig_cgo_3;
  input ensig_cgo_4;



  // Interconnect Declarations for Component Instantiations 
  assign W_tiling_unit_L3_run_cmp_ccs_ccore_en = run_wen & (ensig_cgo | ensig_cgo_iro);
  assign W_tiling_unit_L2_run_cmp_ccs_ccore_en = run_wen & (ensig_cgo_1 | ensig_cgo_iro_1);
  assign O_tiling_unit_L3_run_cmp_ccs_ccore_en = run_wen & (ensig_cgo_2 | ensig_cgo_iro_2);
  assign O_tiling_unit_L2_run_cmp_ccs_ccore_en = run_wen & (ensig_cgo_3 | ensig_cgo_iro_3);
  assign O_tiling_unit_L1_run_cmp_ccs_ccore_en = run_wen & (ensig_cgo_4 | ensig_cgo_iro_4);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci_W_instr_L3_out_wait_dp
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci_W_instr_L3_out_wait_dp
    (
  clk, rst, W_instr_L3_out_rsci_oswt, W_instr_L3_out_rsci_wen_comp, W_instr_L3_out_rsci_biwt,
      W_instr_L3_out_rsci_bdwt, W_instr_L3_out_rsci_bcwt
);
  input clk;
  input rst;
  input W_instr_L3_out_rsci_oswt;
  output W_instr_L3_out_rsci_wen_comp;
  input W_instr_L3_out_rsci_biwt;
  input W_instr_L3_out_rsci_bdwt;
  output W_instr_L3_out_rsci_bcwt;
  reg W_instr_L3_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign W_instr_L3_out_rsci_wen_comp = (~ W_instr_L3_out_rsci_oswt) | W_instr_L3_out_rsci_biwt
      | W_instr_L3_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      W_instr_L3_out_rsci_bcwt <= 1'b0;
    end
    else begin
      W_instr_L3_out_rsci_bcwt <= ~((~(W_instr_L3_out_rsci_bcwt | W_instr_L3_out_rsci_biwt))
          | W_instr_L3_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci_W_instr_L3_out_wait_ctrl
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci_W_instr_L3_out_wait_ctrl
    (
  run_wen, W_instr_L3_out_rsci_oswt, W_instr_L3_out_rsci_irdy, W_instr_L3_out_rsci_biwt,
      W_instr_L3_out_rsci_bdwt, W_instr_L3_out_rsci_bcwt, W_instr_L3_out_rsci_ivld_run_sct
);
  input run_wen;
  input W_instr_L3_out_rsci_oswt;
  input W_instr_L3_out_rsci_irdy;
  output W_instr_L3_out_rsci_biwt;
  output W_instr_L3_out_rsci_bdwt;
  input W_instr_L3_out_rsci_bcwt;
  output W_instr_L3_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire W_instr_L3_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign W_instr_L3_out_rsci_bdwt = W_instr_L3_out_rsci_oswt & run_wen;
  assign W_instr_L3_out_rsci_biwt = W_instr_L3_out_rsci_ogwt & W_instr_L3_out_rsci_irdy;
  assign W_instr_L3_out_rsci_ogwt = W_instr_L3_out_rsci_oswt & (~ W_instr_L3_out_rsci_bcwt);
  assign W_instr_L3_out_rsci_ivld_run_sct = W_instr_L3_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci_W_instr_L2_out_wait_dp
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci_W_instr_L2_out_wait_dp
    (
  clk, rst, W_instr_L2_out_rsci_oswt, W_instr_L2_out_rsci_wen_comp, W_instr_L2_out_rsci_biwt,
      W_instr_L2_out_rsci_bdwt, W_instr_L2_out_rsci_bcwt
);
  input clk;
  input rst;
  input W_instr_L2_out_rsci_oswt;
  output W_instr_L2_out_rsci_wen_comp;
  input W_instr_L2_out_rsci_biwt;
  input W_instr_L2_out_rsci_bdwt;
  output W_instr_L2_out_rsci_bcwt;
  reg W_instr_L2_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign W_instr_L2_out_rsci_wen_comp = (~ W_instr_L2_out_rsci_oswt) | W_instr_L2_out_rsci_biwt
      | W_instr_L2_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      W_instr_L2_out_rsci_bcwt <= 1'b0;
    end
    else begin
      W_instr_L2_out_rsci_bcwt <= ~((~(W_instr_L2_out_rsci_bcwt | W_instr_L2_out_rsci_biwt))
          | W_instr_L2_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci_W_instr_L2_out_wait_ctrl
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci_W_instr_L2_out_wait_ctrl
    (
  run_wen, W_instr_L2_out_rsci_oswt, W_instr_L2_out_rsci_irdy, W_instr_L2_out_rsci_biwt,
      W_instr_L2_out_rsci_bdwt, W_instr_L2_out_rsci_bcwt, W_instr_L2_out_rsci_ivld_run_sct
);
  input run_wen;
  input W_instr_L2_out_rsci_oswt;
  input W_instr_L2_out_rsci_irdy;
  output W_instr_L2_out_rsci_biwt;
  output W_instr_L2_out_rsci_bdwt;
  input W_instr_L2_out_rsci_bcwt;
  output W_instr_L2_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire W_instr_L2_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign W_instr_L2_out_rsci_bdwt = W_instr_L2_out_rsci_oswt & run_wen;
  assign W_instr_L2_out_rsci_biwt = W_instr_L2_out_rsci_ogwt & W_instr_L2_out_rsci_irdy;
  assign W_instr_L2_out_rsci_ogwt = W_instr_L2_out_rsci_oswt & (~ W_instr_L2_out_rsci_bcwt);
  assign W_instr_L2_out_rsci_ivld_run_sct = W_instr_L2_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci_W_instr_L1_out_wait_dp
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci_W_instr_L1_out_wait_dp
    (
  clk, rst, W_instr_L1_out_rsci_oswt, W_instr_L1_out_rsci_wen_comp, W_instr_L1_out_rsci_biwt,
      W_instr_L1_out_rsci_bdwt, W_instr_L1_out_rsci_bcwt
);
  input clk;
  input rst;
  input W_instr_L1_out_rsci_oswt;
  output W_instr_L1_out_rsci_wen_comp;
  input W_instr_L1_out_rsci_biwt;
  input W_instr_L1_out_rsci_bdwt;
  output W_instr_L1_out_rsci_bcwt;
  reg W_instr_L1_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign W_instr_L1_out_rsci_wen_comp = (~ W_instr_L1_out_rsci_oswt) | W_instr_L1_out_rsci_biwt
      | W_instr_L1_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      W_instr_L1_out_rsci_bcwt <= 1'b0;
    end
    else begin
      W_instr_L1_out_rsci_bcwt <= ~((~(W_instr_L1_out_rsci_bcwt | W_instr_L1_out_rsci_biwt))
          | W_instr_L1_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci_W_instr_L1_out_wait_ctrl
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci_W_instr_L1_out_wait_ctrl
    (
  run_wen, W_instr_L1_out_rsci_oswt, W_instr_L1_out_rsci_irdy, W_instr_L1_out_rsci_biwt,
      W_instr_L1_out_rsci_bdwt, W_instr_L1_out_rsci_bcwt, W_instr_L1_out_rsci_ivld_run_sct
);
  input run_wen;
  input W_instr_L1_out_rsci_oswt;
  input W_instr_L1_out_rsci_irdy;
  output W_instr_L1_out_rsci_biwt;
  output W_instr_L1_out_rsci_bdwt;
  input W_instr_L1_out_rsci_bcwt;
  output W_instr_L1_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire W_instr_L1_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign W_instr_L1_out_rsci_bdwt = W_instr_L1_out_rsci_oswt & run_wen;
  assign W_instr_L1_out_rsci_biwt = W_instr_L1_out_rsci_ogwt & W_instr_L1_out_rsci_irdy;
  assign W_instr_L1_out_rsci_ogwt = W_instr_L1_out_rsci_oswt & (~ W_instr_L1_out_rsci_bcwt);
  assign W_instr_L1_out_rsci_ivld_run_sct = W_instr_L1_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci_I_instr_L3_out_wait_dp
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci_I_instr_L3_out_wait_dp
    (
  clk, rst, I_instr_L3_out_rsci_oswt, I_instr_L3_out_rsci_wen_comp, I_instr_L3_out_rsci_biwt,
      I_instr_L3_out_rsci_bdwt, I_instr_L3_out_rsci_bcwt
);
  input clk;
  input rst;
  input I_instr_L3_out_rsci_oswt;
  output I_instr_L3_out_rsci_wen_comp;
  input I_instr_L3_out_rsci_biwt;
  input I_instr_L3_out_rsci_bdwt;
  output I_instr_L3_out_rsci_bcwt;
  reg I_instr_L3_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign I_instr_L3_out_rsci_wen_comp = (~ I_instr_L3_out_rsci_oswt) | I_instr_L3_out_rsci_biwt
      | I_instr_L3_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      I_instr_L3_out_rsci_bcwt <= 1'b0;
    end
    else begin
      I_instr_L3_out_rsci_bcwt <= ~((~(I_instr_L3_out_rsci_bcwt | I_instr_L3_out_rsci_biwt))
          | I_instr_L3_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci_I_instr_L3_out_wait_ctrl
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci_I_instr_L3_out_wait_ctrl
    (
  run_wen, I_instr_L3_out_rsci_oswt, I_instr_L3_out_rsci_irdy, I_instr_L3_out_rsci_biwt,
      I_instr_L3_out_rsci_bdwt, I_instr_L3_out_rsci_bcwt, I_instr_L3_out_rsci_ivld_run_sct
);
  input run_wen;
  input I_instr_L3_out_rsci_oswt;
  input I_instr_L3_out_rsci_irdy;
  output I_instr_L3_out_rsci_biwt;
  output I_instr_L3_out_rsci_bdwt;
  input I_instr_L3_out_rsci_bcwt;
  output I_instr_L3_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire I_instr_L3_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign I_instr_L3_out_rsci_bdwt = I_instr_L3_out_rsci_oswt & run_wen;
  assign I_instr_L3_out_rsci_biwt = I_instr_L3_out_rsci_ogwt & I_instr_L3_out_rsci_irdy;
  assign I_instr_L3_out_rsci_ogwt = I_instr_L3_out_rsci_oswt & (~ I_instr_L3_out_rsci_bcwt);
  assign I_instr_L3_out_rsci_ivld_run_sct = I_instr_L3_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci_I_instr_L2_out_wait_dp
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci_I_instr_L2_out_wait_dp
    (
  clk, rst, I_instr_L2_out_rsci_oswt, I_instr_L2_out_rsci_wen_comp, I_instr_L2_out_rsci_biwt,
      I_instr_L2_out_rsci_bdwt, I_instr_L2_out_rsci_bcwt
);
  input clk;
  input rst;
  input I_instr_L2_out_rsci_oswt;
  output I_instr_L2_out_rsci_wen_comp;
  input I_instr_L2_out_rsci_biwt;
  input I_instr_L2_out_rsci_bdwt;
  output I_instr_L2_out_rsci_bcwt;
  reg I_instr_L2_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign I_instr_L2_out_rsci_wen_comp = (~ I_instr_L2_out_rsci_oswt) | I_instr_L2_out_rsci_biwt
      | I_instr_L2_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      I_instr_L2_out_rsci_bcwt <= 1'b0;
    end
    else begin
      I_instr_L2_out_rsci_bcwt <= ~((~(I_instr_L2_out_rsci_bcwt | I_instr_L2_out_rsci_biwt))
          | I_instr_L2_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci_I_instr_L2_out_wait_ctrl
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci_I_instr_L2_out_wait_ctrl
    (
  run_wen, I_instr_L2_out_rsci_oswt, I_instr_L2_out_rsci_irdy, I_instr_L2_out_rsci_biwt,
      I_instr_L2_out_rsci_bdwt, I_instr_L2_out_rsci_bcwt, I_instr_L2_out_rsci_ivld_run_sct
);
  input run_wen;
  input I_instr_L2_out_rsci_oswt;
  input I_instr_L2_out_rsci_irdy;
  output I_instr_L2_out_rsci_biwt;
  output I_instr_L2_out_rsci_bdwt;
  input I_instr_L2_out_rsci_bcwt;
  output I_instr_L2_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire I_instr_L2_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign I_instr_L2_out_rsci_bdwt = I_instr_L2_out_rsci_oswt & run_wen;
  assign I_instr_L2_out_rsci_biwt = I_instr_L2_out_rsci_ogwt & I_instr_L2_out_rsci_irdy;
  assign I_instr_L2_out_rsci_ogwt = I_instr_L2_out_rsci_oswt & (~ I_instr_L2_out_rsci_bcwt);
  assign I_instr_L2_out_rsci_ivld_run_sct = I_instr_L2_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci_I_instr_L1_out_wait_dp
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci_I_instr_L1_out_wait_dp
    (
  clk, rst, I_instr_L1_out_rsci_oswt, I_instr_L1_out_rsci_wen_comp, I_instr_L1_out_rsci_biwt,
      I_instr_L1_out_rsci_bdwt, I_instr_L1_out_rsci_bcwt
);
  input clk;
  input rst;
  input I_instr_L1_out_rsci_oswt;
  output I_instr_L1_out_rsci_wen_comp;
  input I_instr_L1_out_rsci_biwt;
  input I_instr_L1_out_rsci_bdwt;
  output I_instr_L1_out_rsci_bcwt;
  reg I_instr_L1_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign I_instr_L1_out_rsci_wen_comp = (~ I_instr_L1_out_rsci_oswt) | I_instr_L1_out_rsci_biwt
      | I_instr_L1_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      I_instr_L1_out_rsci_bcwt <= 1'b0;
    end
    else begin
      I_instr_L1_out_rsci_bcwt <= ~((~(I_instr_L1_out_rsci_bcwt | I_instr_L1_out_rsci_biwt))
          | I_instr_L1_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci_I_instr_L1_out_wait_ctrl
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci_I_instr_L1_out_wait_ctrl
    (
  run_wen, I_instr_L1_out_rsci_oswt, I_instr_L1_out_rsci_irdy, I_instr_L1_out_rsci_biwt,
      I_instr_L1_out_rsci_bdwt, I_instr_L1_out_rsci_bcwt, I_instr_L1_out_rsci_ivld_run_sct
);
  input run_wen;
  input I_instr_L1_out_rsci_oswt;
  input I_instr_L1_out_rsci_irdy;
  output I_instr_L1_out_rsci_biwt;
  output I_instr_L1_out_rsci_bdwt;
  input I_instr_L1_out_rsci_bcwt;
  output I_instr_L1_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire I_instr_L1_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign I_instr_L1_out_rsci_bdwt = I_instr_L1_out_rsci_oswt & run_wen;
  assign I_instr_L1_out_rsci_biwt = I_instr_L1_out_rsci_ogwt & I_instr_L1_out_rsci_irdy;
  assign I_instr_L1_out_rsci_ogwt = I_instr_L1_out_rsci_oswt & (~ I_instr_L1_out_rsci_bcwt);
  assign I_instr_L1_out_rsci_ivld_run_sct = I_instr_L1_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci_O_instr_L3_out_wait_dp
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci_O_instr_L3_out_wait_dp
    (
  clk, rst, O_instr_L3_out_rsci_oswt, O_instr_L3_out_rsci_wen_comp, O_instr_L3_out_rsci_biwt,
      O_instr_L3_out_rsci_bdwt, O_instr_L3_out_rsci_bcwt
);
  input clk;
  input rst;
  input O_instr_L3_out_rsci_oswt;
  output O_instr_L3_out_rsci_wen_comp;
  input O_instr_L3_out_rsci_biwt;
  input O_instr_L3_out_rsci_bdwt;
  output O_instr_L3_out_rsci_bcwt;
  reg O_instr_L3_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign O_instr_L3_out_rsci_wen_comp = (~ O_instr_L3_out_rsci_oswt) | O_instr_L3_out_rsci_biwt
      | O_instr_L3_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      O_instr_L3_out_rsci_bcwt <= 1'b0;
    end
    else begin
      O_instr_L3_out_rsci_bcwt <= ~((~(O_instr_L3_out_rsci_bcwt | O_instr_L3_out_rsci_biwt))
          | O_instr_L3_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci_O_instr_L3_out_wait_ctrl
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci_O_instr_L3_out_wait_ctrl
    (
  run_wen, O_instr_L3_out_rsci_oswt, O_instr_L3_out_rsci_irdy, O_instr_L3_out_rsci_biwt,
      O_instr_L3_out_rsci_bdwt, O_instr_L3_out_rsci_bcwt, O_instr_L3_out_rsci_ivld_run_sct
);
  input run_wen;
  input O_instr_L3_out_rsci_oswt;
  input O_instr_L3_out_rsci_irdy;
  output O_instr_L3_out_rsci_biwt;
  output O_instr_L3_out_rsci_bdwt;
  input O_instr_L3_out_rsci_bcwt;
  output O_instr_L3_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire O_instr_L3_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign O_instr_L3_out_rsci_bdwt = O_instr_L3_out_rsci_oswt & run_wen;
  assign O_instr_L3_out_rsci_biwt = O_instr_L3_out_rsci_ogwt & O_instr_L3_out_rsci_irdy;
  assign O_instr_L3_out_rsci_ogwt = O_instr_L3_out_rsci_oswt & (~ O_instr_L3_out_rsci_bcwt);
  assign O_instr_L3_out_rsci_ivld_run_sct = O_instr_L3_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci_O_instr_L2_out_wait_dp
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci_O_instr_L2_out_wait_dp
    (
  clk, rst, O_instr_L2_out_rsci_oswt, O_instr_L2_out_rsci_wen_comp, O_instr_L2_out_rsci_biwt,
      O_instr_L2_out_rsci_bdwt, O_instr_L2_out_rsci_bcwt
);
  input clk;
  input rst;
  input O_instr_L2_out_rsci_oswt;
  output O_instr_L2_out_rsci_wen_comp;
  input O_instr_L2_out_rsci_biwt;
  input O_instr_L2_out_rsci_bdwt;
  output O_instr_L2_out_rsci_bcwt;
  reg O_instr_L2_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign O_instr_L2_out_rsci_wen_comp = (~ O_instr_L2_out_rsci_oswt) | O_instr_L2_out_rsci_biwt
      | O_instr_L2_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      O_instr_L2_out_rsci_bcwt <= 1'b0;
    end
    else begin
      O_instr_L2_out_rsci_bcwt <= ~((~(O_instr_L2_out_rsci_bcwt | O_instr_L2_out_rsci_biwt))
          | O_instr_L2_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci_O_instr_L2_out_wait_ctrl
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci_O_instr_L2_out_wait_ctrl
    (
  run_wen, O_instr_L2_out_rsci_oswt, O_instr_L2_out_rsci_irdy, O_instr_L2_out_rsci_biwt,
      O_instr_L2_out_rsci_bdwt, O_instr_L2_out_rsci_bcwt, O_instr_L2_out_rsci_ivld_run_sct
);
  input run_wen;
  input O_instr_L2_out_rsci_oswt;
  input O_instr_L2_out_rsci_irdy;
  output O_instr_L2_out_rsci_biwt;
  output O_instr_L2_out_rsci_bdwt;
  input O_instr_L2_out_rsci_bcwt;
  output O_instr_L2_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire O_instr_L2_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign O_instr_L2_out_rsci_bdwt = O_instr_L2_out_rsci_oswt & run_wen;
  assign O_instr_L2_out_rsci_biwt = O_instr_L2_out_rsci_ogwt & O_instr_L2_out_rsci_irdy;
  assign O_instr_L2_out_rsci_ogwt = O_instr_L2_out_rsci_oswt & (~ O_instr_L2_out_rsci_bcwt);
  assign O_instr_L2_out_rsci_ivld_run_sct = O_instr_L2_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci_O_instr_L1_out_wait_dp
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci_O_instr_L1_out_wait_dp
    (
  clk, rst, O_instr_L1_out_rsci_oswt, O_instr_L1_out_rsci_wen_comp, O_instr_L1_out_rsci_biwt,
      O_instr_L1_out_rsci_bdwt, O_instr_L1_out_rsci_bcwt
);
  input clk;
  input rst;
  input O_instr_L1_out_rsci_oswt;
  output O_instr_L1_out_rsci_wen_comp;
  input O_instr_L1_out_rsci_biwt;
  input O_instr_L1_out_rsci_bdwt;
  output O_instr_L1_out_rsci_bcwt;
  reg O_instr_L1_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign O_instr_L1_out_rsci_wen_comp = (~ O_instr_L1_out_rsci_oswt) | O_instr_L1_out_rsci_biwt
      | O_instr_L1_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      O_instr_L1_out_rsci_bcwt <= 1'b0;
    end
    else begin
      O_instr_L1_out_rsci_bcwt <= ~((~(O_instr_L1_out_rsci_bcwt | O_instr_L1_out_rsci_biwt))
          | O_instr_L1_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci_O_instr_L1_out_wait_ctrl
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci_O_instr_L1_out_wait_ctrl
    (
  run_wen, O_instr_L1_out_rsci_oswt, O_instr_L1_out_rsci_irdy, O_instr_L1_out_rsci_biwt,
      O_instr_L1_out_rsci_bdwt, O_instr_L1_out_rsci_bcwt, O_instr_L1_out_rsci_ivld_run_sct
);
  input run_wen;
  input O_instr_L1_out_rsci_oswt;
  input O_instr_L1_out_rsci_irdy;
  output O_instr_L1_out_rsci_biwt;
  output O_instr_L1_out_rsci_bdwt;
  input O_instr_L1_out_rsci_bcwt;
  output O_instr_L1_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire O_instr_L1_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign O_instr_L1_out_rsci_bdwt = O_instr_L1_out_rsci_oswt & run_wen;
  assign O_instr_L1_out_rsci_biwt = O_instr_L1_out_rsci_ogwt & O_instr_L1_out_rsci_irdy;
  assign O_instr_L1_out_rsci_ogwt = O_instr_L1_out_rsci_oswt & (~ O_instr_L1_out_rsci_bcwt);
  assign O_instr_L1_out_rsci_ivld_run_sct = O_instr_L1_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_layer_instruction_in_rsci_layer_instruction_in_wait_dp
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_layer_instruction_in_rsci_layer_instruction_in_wait_dp
    (
  clk, rst, layer_instruction_in_rsci_oswt, layer_instruction_in_rsci_wen_comp, layer_instruction_in_rsci_idat_mxwt,
      layer_instruction_in_rsci_biwt, layer_instruction_in_rsci_bdwt, layer_instruction_in_rsci_bcwt,
      layer_instruction_in_rsci_idat
);
  input clk;
  input rst;
  input layer_instruction_in_rsci_oswt;
  output layer_instruction_in_rsci_wen_comp;
  output [484:0] layer_instruction_in_rsci_idat_mxwt;
  input layer_instruction_in_rsci_biwt;
  input layer_instruction_in_rsci_bdwt;
  output layer_instruction_in_rsci_bcwt;
  reg layer_instruction_in_rsci_bcwt;
  input [484:0] layer_instruction_in_rsci_idat;


  // Interconnect Declarations
  reg [484:0] layer_instruction_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign layer_instruction_in_rsci_wen_comp = (~ layer_instruction_in_rsci_oswt)
      | layer_instruction_in_rsci_biwt | layer_instruction_in_rsci_bcwt;
  assign layer_instruction_in_rsci_idat_mxwt = MUX_v_485_2_2(layer_instruction_in_rsci_idat,
      layer_instruction_in_rsci_idat_bfwt, layer_instruction_in_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      layer_instruction_in_rsci_bcwt <= 1'b0;
    end
    else begin
      layer_instruction_in_rsci_bcwt <= ~((~(layer_instruction_in_rsci_bcwt | layer_instruction_in_rsci_biwt))
          | layer_instruction_in_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer_instruction_in_rsci_idat_bfwt <= 485'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( layer_instruction_in_rsci_biwt ) begin
      layer_instruction_in_rsci_idat_bfwt <= layer_instruction_in_rsci_idat;
    end
  end

  function automatic [484:0] MUX_v_485_2_2;
    input [484:0] input_0;
    input [484:0] input_1;
    input [0:0] sel;
    reg [484:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_485_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_layer_instruction_in_rsci_layer_instruction_in_wait_ctrl
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_layer_instruction_in_rsci_layer_instruction_in_wait_ctrl
    (
  run_wen, layer_instruction_in_rsci_oswt, layer_instruction_in_rsci_biwt, layer_instruction_in_rsci_bdwt,
      layer_instruction_in_rsci_bcwt, layer_instruction_in_rsci_irdy_run_sct, layer_instruction_in_rsci_ivld
);
  input run_wen;
  input layer_instruction_in_rsci_oswt;
  output layer_instruction_in_rsci_biwt;
  output layer_instruction_in_rsci_bdwt;
  input layer_instruction_in_rsci_bcwt;
  output layer_instruction_in_rsci_irdy_run_sct;
  input layer_instruction_in_rsci_ivld;


  // Interconnect Declarations
  wire layer_instruction_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign layer_instruction_in_rsci_bdwt = layer_instruction_in_rsci_oswt & run_wen;
  assign layer_instruction_in_rsci_biwt = layer_instruction_in_rsci_ogwt & layer_instruction_in_rsci_ivld;
  assign layer_instruction_in_rsci_ogwt = layer_instruction_in_rsci_oswt & (~ layer_instruction_in_rsci_bcwt);
  assign layer_instruction_in_rsci_irdy_run_sct = layer_instruction_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_run_fsm
    (
  clk, rst, run_wen, fsm_output
);
  input clk;
  input rst;
  input run_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_run_fsm_1
  parameter
    run_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_staller
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_staller
    (
  clk, rst, run_wen, run_wten, O_instr_in_rsci_wen_comp, I_instr_in_rsci_wen_comp,
      W_instr_in_rsci_wen_comp
);
  input clk;
  input rst;
  output run_wen;
  output run_wten;
  reg run_wten;
  input O_instr_in_rsci_wen_comp;
  input I_instr_in_rsci_wen_comp;
  input W_instr_in_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = O_instr_in_rsci_wen_comp & I_instr_in_rsci_wen_comp & W_instr_in_rsci_wen_comp;
  always @(posedge clk) begin
    if ( rst ) begin
      run_wten <= 1'b0;
    end
    else begin
      run_wten <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_instr_in_rsci_W_instr_in_wait_dp
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_instr_in_rsci_W_instr_in_wait_dp
    (
  clk, rst, W_instr_in_rsci_oswt, W_instr_in_rsci_wen_comp, W_instr_in_rsci_idat_mxwt,
      W_instr_in_rsci_biwt, W_instr_in_rsci_bdwt, W_instr_in_rsci_bcwt, W_instr_in_rsci_idat
);
  input clk;
  input rst;
  input W_instr_in_rsci_oswt;
  output W_instr_in_rsci_wen_comp;
  output [49:0] W_instr_in_rsci_idat_mxwt;
  input W_instr_in_rsci_biwt;
  input W_instr_in_rsci_bdwt;
  output W_instr_in_rsci_bcwt;
  reg W_instr_in_rsci_bcwt;
  input [49:0] W_instr_in_rsci_idat;


  // Interconnect Declarations
  reg [49:0] W_instr_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign W_instr_in_rsci_wen_comp = (~ W_instr_in_rsci_oswt) | W_instr_in_rsci_biwt
      | W_instr_in_rsci_bcwt;
  assign W_instr_in_rsci_idat_mxwt = MUX_v_50_2_2(W_instr_in_rsci_idat, W_instr_in_rsci_idat_bfwt,
      W_instr_in_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      W_instr_in_rsci_bcwt <= 1'b0;
    end
    else begin
      W_instr_in_rsci_bcwt <= ~((~(W_instr_in_rsci_bcwt | W_instr_in_rsci_biwt))
          | W_instr_in_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_instr_in_rsci_idat_bfwt <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( W_instr_in_rsci_biwt ) begin
      W_instr_in_rsci_idat_bfwt <= W_instr_in_rsci_idat;
    end
  end

  function automatic [49:0] MUX_v_50_2_2;
    input [49:0] input_0;
    input [49:0] input_1;
    input [0:0] sel;
    reg [49:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_50_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_instr_in_rsci_W_instr_in_wait_ctrl
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_instr_in_rsci_W_instr_in_wait_ctrl
    (
  run_wen, W_instr_in_rsci_oswt, W_instr_in_rsci_biwt, W_instr_in_rsci_bdwt, W_instr_in_rsci_bcwt,
      W_instr_in_rsci_irdy_run_sct, W_instr_in_rsci_ivld
);
  input run_wen;
  input W_instr_in_rsci_oswt;
  output W_instr_in_rsci_biwt;
  output W_instr_in_rsci_bdwt;
  input W_instr_in_rsci_bcwt;
  output W_instr_in_rsci_irdy_run_sct;
  input W_instr_in_rsci_ivld;


  // Interconnect Declarations
  wire W_instr_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign W_instr_in_rsci_bdwt = W_instr_in_rsci_oswt & run_wen;
  assign W_instr_in_rsci_biwt = W_instr_in_rsci_ogwt & W_instr_in_rsci_ivld;
  assign W_instr_in_rsci_ogwt = W_instr_in_rsci_oswt & (~ W_instr_in_rsci_bcwt);
  assign W_instr_in_rsci_irdy_run_sct = W_instr_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_instr_in_rsci_I_instr_in_wait_dp
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_instr_in_rsci_I_instr_in_wait_dp
    (
  clk, rst, I_instr_in_rsci_oswt, I_instr_in_rsci_wen_comp, I_instr_in_rsci_idat_mxwt,
      I_instr_in_rsci_biwt, I_instr_in_rsci_bdwt, I_instr_in_rsci_bcwt, I_instr_in_rsci_idat
);
  input clk;
  input rst;
  input I_instr_in_rsci_oswt;
  output I_instr_in_rsci_wen_comp;
  output [49:0] I_instr_in_rsci_idat_mxwt;
  input I_instr_in_rsci_biwt;
  input I_instr_in_rsci_bdwt;
  output I_instr_in_rsci_bcwt;
  reg I_instr_in_rsci_bcwt;
  input [49:0] I_instr_in_rsci_idat;


  // Interconnect Declarations
  reg [49:0] I_instr_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign I_instr_in_rsci_wen_comp = (~ I_instr_in_rsci_oswt) | I_instr_in_rsci_biwt
      | I_instr_in_rsci_bcwt;
  assign I_instr_in_rsci_idat_mxwt = MUX_v_50_2_2(I_instr_in_rsci_idat, I_instr_in_rsci_idat_bfwt,
      I_instr_in_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      I_instr_in_rsci_bcwt <= 1'b0;
    end
    else begin
      I_instr_in_rsci_bcwt <= ~((~(I_instr_in_rsci_bcwt | I_instr_in_rsci_biwt))
          | I_instr_in_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_instr_in_rsci_idat_bfwt <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( I_instr_in_rsci_biwt ) begin
      I_instr_in_rsci_idat_bfwt <= I_instr_in_rsci_idat;
    end
  end

  function automatic [49:0] MUX_v_50_2_2;
    input [49:0] input_0;
    input [49:0] input_1;
    input [0:0] sel;
    reg [49:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_50_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_instr_in_rsci_I_instr_in_wait_ctrl
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_instr_in_rsci_I_instr_in_wait_ctrl
    (
  run_wen, I_instr_in_rsci_oswt, I_instr_in_rsci_biwt, I_instr_in_rsci_bdwt, I_instr_in_rsci_bcwt,
      I_instr_in_rsci_irdy_run_sct, I_instr_in_rsci_ivld
);
  input run_wen;
  input I_instr_in_rsci_oswt;
  output I_instr_in_rsci_biwt;
  output I_instr_in_rsci_bdwt;
  input I_instr_in_rsci_bcwt;
  output I_instr_in_rsci_irdy_run_sct;
  input I_instr_in_rsci_ivld;


  // Interconnect Declarations
  wire I_instr_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign I_instr_in_rsci_bdwt = I_instr_in_rsci_oswt & run_wen;
  assign I_instr_in_rsci_biwt = I_instr_in_rsci_ogwt & I_instr_in_rsci_ivld;
  assign I_instr_in_rsci_ogwt = I_instr_in_rsci_oswt & (~ I_instr_in_rsci_bcwt);
  assign I_instr_in_rsci_irdy_run_sct = I_instr_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_instr_in_rsci_O_instr_in_wait_dp
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_instr_in_rsci_O_instr_in_wait_dp
    (
  clk, rst, O_instr_in_rsci_oswt, O_instr_in_rsci_wen_comp, O_instr_in_rsci_idat_mxwt,
      O_instr_in_rsci_biwt, O_instr_in_rsci_bdwt, O_instr_in_rsci_bcwt, O_instr_in_rsci_idat
);
  input clk;
  input rst;
  input O_instr_in_rsci_oswt;
  output O_instr_in_rsci_wen_comp;
  output [49:0] O_instr_in_rsci_idat_mxwt;
  input O_instr_in_rsci_biwt;
  input O_instr_in_rsci_bdwt;
  output O_instr_in_rsci_bcwt;
  reg O_instr_in_rsci_bcwt;
  input [49:0] O_instr_in_rsci_idat;


  // Interconnect Declarations
  reg [49:0] O_instr_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign O_instr_in_rsci_wen_comp = (~ O_instr_in_rsci_oswt) | O_instr_in_rsci_biwt
      | O_instr_in_rsci_bcwt;
  assign O_instr_in_rsci_idat_mxwt = MUX_v_50_2_2(O_instr_in_rsci_idat, O_instr_in_rsci_idat_bfwt,
      O_instr_in_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      O_instr_in_rsci_bcwt <= 1'b0;
    end
    else begin
      O_instr_in_rsci_bcwt <= ~((~(O_instr_in_rsci_bcwt | O_instr_in_rsci_biwt))
          | O_instr_in_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_instr_in_rsci_idat_bfwt <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( O_instr_in_rsci_biwt ) begin
      O_instr_in_rsci_idat_bfwt <= O_instr_in_rsci_idat;
    end
  end

  function automatic [49:0] MUX_v_50_2_2;
    input [49:0] input_0;
    input [49:0] input_1;
    input [0:0] sel;
    reg [49:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_50_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_instr_in_rsci_O_instr_in_wait_ctrl
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_instr_in_rsci_O_instr_in_wait_ctrl
    (
  run_wen, O_instr_in_rsci_oswt, O_instr_in_rsci_biwt, O_instr_in_rsci_bdwt, O_instr_in_rsci_bcwt,
      O_instr_in_rsci_irdy_run_sct, O_instr_in_rsci_ivld
);
  input run_wen;
  input O_instr_in_rsci_oswt;
  output O_instr_in_rsci_biwt;
  output O_instr_in_rsci_bdwt;
  input O_instr_in_rsci_bcwt;
  output O_instr_in_rsci_irdy_run_sct;
  input O_instr_in_rsci_ivld;


  // Interconnect Declarations
  wire O_instr_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign O_instr_in_rsci_bdwt = O_instr_in_rsci_oswt & run_wen;
  assign O_instr_in_rsci_biwt = O_instr_in_rsci_ogwt & O_instr_in_rsci_ivld;
  assign O_instr_in_rsci_ogwt = O_instr_in_rsci_oswt & (~ O_instr_in_rsci_bcwt);
  assign O_instr_in_rsci_irdy_run_sct = O_instr_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_wr_data_zero_guard_rsci_wr_data_zero_guard_wait_dp
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_wr_data_zero_guard_rsci_wr_data_zero_guard_wait_dp
    (
  clk, rst, wr_data_zero_guard_rsci_ivld_mxwt, wr_data_zero_guard_rsci_idat_mxwt,
      wr_data_zero_guard_rsci_biwt, wr_data_zero_guard_rsci_bdwt, wr_data_zero_guard_rsci_ivld,
      wr_data_zero_guard_rsci_idat
);
  input clk;
  input rst;
  output wr_data_zero_guard_rsci_ivld_mxwt;
  output wr_data_zero_guard_rsci_idat_mxwt;
  input wr_data_zero_guard_rsci_biwt;
  input wr_data_zero_guard_rsci_bdwt;
  input wr_data_zero_guard_rsci_ivld;
  input wr_data_zero_guard_rsci_idat;


  // Interconnect Declarations
  reg wr_data_zero_guard_rsci_bcwt;
  reg wr_data_zero_guard_rsci_ivld_bfwt;
  wire wr_data_zero_guard_rsci_idat_gtd;
  reg wr_data_zero_guard_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign wr_data_zero_guard_rsci_ivld_mxwt = MUX_s_1_2_2(wr_data_zero_guard_rsci_ivld,
      wr_data_zero_guard_rsci_ivld_bfwt, wr_data_zero_guard_rsci_bcwt);
  assign wr_data_zero_guard_rsci_idat_gtd = wr_data_zero_guard_rsci_idat & wr_data_zero_guard_rsci_ivld;
  assign wr_data_zero_guard_rsci_idat_mxwt = MUX_s_1_2_2(wr_data_zero_guard_rsci_idat_gtd,
      wr_data_zero_guard_rsci_idat_bfwt, wr_data_zero_guard_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      wr_data_zero_guard_rsci_bcwt <= 1'b0;
    end
    else begin
      wr_data_zero_guard_rsci_bcwt <= ~((~(wr_data_zero_guard_rsci_bcwt | wr_data_zero_guard_rsci_biwt))
          | wr_data_zero_guard_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      wr_data_zero_guard_rsci_ivld_bfwt <= 1'b0;
      wr_data_zero_guard_rsci_idat_bfwt <= 1'b0;
    end
    else if ( wr_data_zero_guard_rsci_biwt ) begin
      wr_data_zero_guard_rsci_ivld_bfwt <= wr_data_zero_guard_rsci_ivld;
      wr_data_zero_guard_rsci_idat_bfwt <= wr_data_zero_guard_rsci_idat_gtd;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_wr_data_zero_guard_rsci_wr_data_zero_guard_wait_ctrl
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_wr_data_zero_guard_rsci_wr_data_zero_guard_wait_ctrl
    (
  run_wen, run_wten, wr_data_zero_guard_rsci_oswt, wr_data_zero_guard_rsci_biwt,
      wr_data_zero_guard_rsci_bdwt
);
  input run_wen;
  input run_wten;
  input wr_data_zero_guard_rsci_oswt;
  output wr_data_zero_guard_rsci_biwt;
  output wr_data_zero_guard_rsci_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign wr_data_zero_guard_rsci_bdwt = wr_data_zero_guard_rsci_oswt & run_wen;
  assign wr_data_zero_guard_rsci_biwt = (~ run_wten) & wr_data_zero_guard_rsci_oswt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_wr_data_rsci_W_wr_data_wait_dp
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_wr_data_rsci_W_wr_data_wait_dp
    (
  clk, rst, W_wr_data_rsci_ivld_mxwt, W_wr_data_rsci_idat_mxwt, W_wr_data_rsci_biwt,
      W_wr_data_rsci_bdwt, W_wr_data_rsci_ivld, W_wr_data_rsci_idat
);
  input clk;
  input rst;
  output W_wr_data_rsci_ivld_mxwt;
  output [15:0] W_wr_data_rsci_idat_mxwt;
  input W_wr_data_rsci_biwt;
  input W_wr_data_rsci_bdwt;
  input W_wr_data_rsci_ivld;
  input [15:0] W_wr_data_rsci_idat;


  // Interconnect Declarations
  reg W_wr_data_rsci_bcwt;
  reg W_wr_data_rsci_ivld_bfwt;
  wire [15:0] W_wr_data_rsci_idat_gtd;
  reg [15:0] W_wr_data_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign W_wr_data_rsci_ivld_mxwt = MUX_s_1_2_2(W_wr_data_rsci_ivld, W_wr_data_rsci_ivld_bfwt,
      W_wr_data_rsci_bcwt);
  assign W_wr_data_rsci_idat_gtd = MUX_v_16_2_2(16'b0000000000000000, W_wr_data_rsci_idat,
      W_wr_data_rsci_ivld);
  assign W_wr_data_rsci_idat_mxwt = MUX_v_16_2_2(W_wr_data_rsci_idat_gtd, W_wr_data_rsci_idat_bfwt,
      W_wr_data_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      W_wr_data_rsci_bcwt <= 1'b0;
    end
    else begin
      W_wr_data_rsci_bcwt <= ~((~(W_wr_data_rsci_bcwt | W_wr_data_rsci_biwt)) | W_wr_data_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_wr_data_rsci_ivld_bfwt <= 1'b0;
      W_wr_data_rsci_idat_bfwt <= 16'b0000000000000000;
    end
    else if ( W_wr_data_rsci_biwt ) begin
      W_wr_data_rsci_ivld_bfwt <= W_wr_data_rsci_ivld;
      W_wr_data_rsci_idat_bfwt <= W_wr_data_rsci_idat_gtd;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_wr_data_rsci_W_wr_data_wait_ctrl
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_wr_data_rsci_W_wr_data_wait_ctrl
    (
  run_wen, run_wten, W_wr_data_rsci_oswt, W_wr_data_rsci_biwt, W_wr_data_rsci_bdwt
);
  input run_wen;
  input run_wten;
  input W_wr_data_rsci_oswt;
  output W_wr_data_rsci_biwt;
  output W_wr_data_rsci_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign W_wr_data_rsci_bdwt = W_wr_data_rsci_oswt & run_wen;
  assign W_wr_data_rsci_biwt = (~ run_wten) & W_wr_data_rsci_oswt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_wr_data_rsci_I_wr_data_wait_dp
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_wr_data_rsci_I_wr_data_wait_dp
    (
  clk, rst, I_wr_data_rsci_ivld_mxwt, I_wr_data_rsci_idat_mxwt, I_wr_data_rsci_biwt,
      I_wr_data_rsci_bdwt, I_wr_data_rsci_ivld, I_wr_data_rsci_idat
);
  input clk;
  input rst;
  output I_wr_data_rsci_ivld_mxwt;
  output [15:0] I_wr_data_rsci_idat_mxwt;
  input I_wr_data_rsci_biwt;
  input I_wr_data_rsci_bdwt;
  input I_wr_data_rsci_ivld;
  input [15:0] I_wr_data_rsci_idat;


  // Interconnect Declarations
  reg I_wr_data_rsci_bcwt;
  reg I_wr_data_rsci_ivld_bfwt;
  wire [15:0] I_wr_data_rsci_idat_gtd;
  reg [15:0] I_wr_data_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign I_wr_data_rsci_ivld_mxwt = MUX_s_1_2_2(I_wr_data_rsci_ivld, I_wr_data_rsci_ivld_bfwt,
      I_wr_data_rsci_bcwt);
  assign I_wr_data_rsci_idat_gtd = MUX_v_16_2_2(16'b0000000000000000, I_wr_data_rsci_idat,
      I_wr_data_rsci_ivld);
  assign I_wr_data_rsci_idat_mxwt = MUX_v_16_2_2(I_wr_data_rsci_idat_gtd, I_wr_data_rsci_idat_bfwt,
      I_wr_data_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      I_wr_data_rsci_bcwt <= 1'b0;
    end
    else begin
      I_wr_data_rsci_bcwt <= ~((~(I_wr_data_rsci_bcwt | I_wr_data_rsci_biwt)) | I_wr_data_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_wr_data_rsci_ivld_bfwt <= 1'b0;
      I_wr_data_rsci_idat_bfwt <= 16'b0000000000000000;
    end
    else if ( I_wr_data_rsci_biwt ) begin
      I_wr_data_rsci_ivld_bfwt <= I_wr_data_rsci_ivld;
      I_wr_data_rsci_idat_bfwt <= I_wr_data_rsci_idat_gtd;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_wr_data_rsci_I_wr_data_wait_ctrl
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_wr_data_rsci_I_wr_data_wait_ctrl
    (
  run_wen, run_wten, I_wr_data_rsci_oswt, I_wr_data_rsci_biwt, I_wr_data_rsci_bdwt
);
  input run_wen;
  input run_wten;
  input I_wr_data_rsci_oswt;
  output I_wr_data_rsci_biwt;
  output I_wr_data_rsci_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign I_wr_data_rsci_bdwt = I_wr_data_rsci_oswt & run_wen;
  assign I_wr_data_rsci_biwt = (~ run_wten) & I_wr_data_rsci_oswt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_rd_data_rsci_O_rd_data_wait_dp
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_rd_data_rsci_O_rd_data_wait_dp
    (
  clk, rst, O_rd_data_rsci_irdy_mxwt, O_rd_data_rsci_irdy, O_rd_data_rsci_biwt, O_rd_data_rsci_bdwt
);
  input clk;
  input rst;
  output O_rd_data_rsci_irdy_mxwt;
  input O_rd_data_rsci_irdy;
  input O_rd_data_rsci_biwt;
  input O_rd_data_rsci_bdwt;


  // Interconnect Declarations
  reg O_rd_data_rsci_bcwt;
  reg O_rd_data_rsci_irdy_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign O_rd_data_rsci_irdy_mxwt = MUX_s_1_2_2(O_rd_data_rsci_irdy, O_rd_data_rsci_irdy_bfwt,
      O_rd_data_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      O_rd_data_rsci_bcwt <= 1'b0;
    end
    else begin
      O_rd_data_rsci_bcwt <= ~((~(O_rd_data_rsci_bcwt | O_rd_data_rsci_biwt)) | O_rd_data_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_rd_data_rsci_irdy_bfwt <= 1'b0;
    end
    else if ( O_rd_data_rsci_biwt ) begin
      O_rd_data_rsci_irdy_bfwt <= O_rd_data_rsci_irdy;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_rd_data_rsci_O_rd_data_wait_ctrl
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_rd_data_rsci_O_rd_data_wait_ctrl
    (
  run_wen, run_wten, O_rd_data_rsci_oswt, O_rd_data_rsci_biwt, O_rd_data_rsci_bdwt
);
  input run_wen;
  input run_wten;
  input O_rd_data_rsci_oswt;
  output O_rd_data_rsci_biwt;
  output O_rd_data_rsci_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign O_rd_data_rsci_bdwt = O_rd_data_rsci_oswt & run_wen;
  assign O_rd_data_rsci_biwt = (~ run_wten) & O_rd_data_rsci_oswt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_wr_data_rsci_O_wr_data_wait_dp
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_wr_data_rsci_O_wr_data_wait_dp
    (
  clk, rst, O_wr_data_rsci_ivld_mxwt, O_wr_data_rsci_idat_mxwt, O_wr_data_rsci_biwt,
      O_wr_data_rsci_bdwt, O_wr_data_rsci_ivld, O_wr_data_rsci_idat
);
  input clk;
  input rst;
  output O_wr_data_rsci_ivld_mxwt;
  output [15:0] O_wr_data_rsci_idat_mxwt;
  input O_wr_data_rsci_biwt;
  input O_wr_data_rsci_bdwt;
  input O_wr_data_rsci_ivld;
  input [15:0] O_wr_data_rsci_idat;


  // Interconnect Declarations
  reg O_wr_data_rsci_bcwt;
  reg O_wr_data_rsci_ivld_bfwt;
  wire [15:0] O_wr_data_rsci_idat_gtd;
  reg [15:0] O_wr_data_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign O_wr_data_rsci_ivld_mxwt = MUX_s_1_2_2(O_wr_data_rsci_ivld, O_wr_data_rsci_ivld_bfwt,
      O_wr_data_rsci_bcwt);
  assign O_wr_data_rsci_idat_gtd = MUX_v_16_2_2(16'b0000000000000000, O_wr_data_rsci_idat,
      O_wr_data_rsci_ivld);
  assign O_wr_data_rsci_idat_mxwt = MUX_v_16_2_2(O_wr_data_rsci_idat_gtd, O_wr_data_rsci_idat_bfwt,
      O_wr_data_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      O_wr_data_rsci_bcwt <= 1'b0;
    end
    else begin
      O_wr_data_rsci_bcwt <= ~((~(O_wr_data_rsci_bcwt | O_wr_data_rsci_biwt)) | O_wr_data_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_wr_data_rsci_ivld_bfwt <= 1'b0;
      O_wr_data_rsci_idat_bfwt <= 16'b0000000000000000;
    end
    else if ( O_wr_data_rsci_biwt ) begin
      O_wr_data_rsci_ivld_bfwt <= O_wr_data_rsci_ivld;
      O_wr_data_rsci_idat_bfwt <= O_wr_data_rsci_idat_gtd;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_wr_data_rsci_O_wr_data_wait_ctrl
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_wr_data_rsci_O_wr_data_wait_ctrl
    (
  run_wen, O_wr_data_rsci_oswt, run_wten, O_wr_data_rsci_biwt, O_wr_data_rsci_bdwt
);
  input run_wen;
  input O_wr_data_rsci_oswt;
  input run_wten;
  output O_wr_data_rsci_biwt;
  output O_wr_data_rsci_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign O_wr_data_rsci_bdwt = O_wr_data_rsci_oswt & run_wen;
  assign O_wr_data_rsci_biwt = (~ run_wten) & O_wr_data_rsci_oswt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci
    (
  clk, rst, W_instr_L3_out_rsc_dat, W_instr_L3_out_rsc_vld, W_instr_L3_out_rsc_rdy,
      run_wen, W_instr_L3_out_rsci_oswt, W_instr_L3_out_rsci_wen_comp, W_instr_L3_out_rsci_idat
);
  input clk;
  input rst;
  output [159:0] W_instr_L3_out_rsc_dat;
  output W_instr_L3_out_rsc_vld;
  input W_instr_L3_out_rsc_rdy;
  input run_wen;
  input W_instr_L3_out_rsci_oswt;
  output W_instr_L3_out_rsci_wen_comp;
  input [159:0] W_instr_L3_out_rsci_idat;


  // Interconnect Declarations
  wire W_instr_L3_out_rsci_irdy;
  wire W_instr_L3_out_rsci_biwt;
  wire W_instr_L3_out_rsci_bdwt;
  wire W_instr_L3_out_rsci_bcwt;
  wire W_instr_L3_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd35),
  .width(32'sd160)) W_instr_L3_out_rsci (
      .irdy(W_instr_L3_out_rsci_irdy),
      .ivld(W_instr_L3_out_rsci_ivld_run_sct),
      .idat(W_instr_L3_out_rsci_idat),
      .rdy(W_instr_L3_out_rsc_rdy),
      .vld(W_instr_L3_out_rsc_vld),
      .dat(W_instr_L3_out_rsc_dat)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci_W_instr_L3_out_wait_ctrl
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci_W_instr_L3_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .W_instr_L3_out_rsci_oswt(W_instr_L3_out_rsci_oswt),
      .W_instr_L3_out_rsci_irdy(W_instr_L3_out_rsci_irdy),
      .W_instr_L3_out_rsci_biwt(W_instr_L3_out_rsci_biwt),
      .W_instr_L3_out_rsci_bdwt(W_instr_L3_out_rsci_bdwt),
      .W_instr_L3_out_rsci_bcwt(W_instr_L3_out_rsci_bcwt),
      .W_instr_L3_out_rsci_ivld_run_sct(W_instr_L3_out_rsci_ivld_run_sct)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci_W_instr_L3_out_wait_dp
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci_W_instr_L3_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .W_instr_L3_out_rsci_oswt(W_instr_L3_out_rsci_oswt),
      .W_instr_L3_out_rsci_wen_comp(W_instr_L3_out_rsci_wen_comp),
      .W_instr_L3_out_rsci_biwt(W_instr_L3_out_rsci_biwt),
      .W_instr_L3_out_rsci_bdwt(W_instr_L3_out_rsci_bdwt),
      .W_instr_L3_out_rsci_bcwt(W_instr_L3_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci
    (
  clk, rst, W_instr_L2_out_rsc_dat, W_instr_L2_out_rsc_vld, W_instr_L2_out_rsc_rdy,
      run_wen, W_instr_L2_out_rsci_oswt, W_instr_L2_out_rsci_wen_comp, W_instr_L2_out_rsci_idat
);
  input clk;
  input rst;
  output [109:0] W_instr_L2_out_rsc_dat;
  output W_instr_L2_out_rsc_vld;
  input W_instr_L2_out_rsc_rdy;
  input run_wen;
  input W_instr_L2_out_rsci_oswt;
  output W_instr_L2_out_rsci_wen_comp;
  input [109:0] W_instr_L2_out_rsci_idat;


  // Interconnect Declarations
  wire W_instr_L2_out_rsci_irdy;
  wire W_instr_L2_out_rsci_biwt;
  wire W_instr_L2_out_rsci_bdwt;
  wire W_instr_L2_out_rsci_bcwt;
  wire W_instr_L2_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd34),
  .width(32'sd110)) W_instr_L2_out_rsci (
      .irdy(W_instr_L2_out_rsci_irdy),
      .ivld(W_instr_L2_out_rsci_ivld_run_sct),
      .idat(W_instr_L2_out_rsci_idat),
      .rdy(W_instr_L2_out_rsc_rdy),
      .vld(W_instr_L2_out_rsc_vld),
      .dat(W_instr_L2_out_rsc_dat)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci_W_instr_L2_out_wait_ctrl
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci_W_instr_L2_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .W_instr_L2_out_rsci_oswt(W_instr_L2_out_rsci_oswt),
      .W_instr_L2_out_rsci_irdy(W_instr_L2_out_rsci_irdy),
      .W_instr_L2_out_rsci_biwt(W_instr_L2_out_rsci_biwt),
      .W_instr_L2_out_rsci_bdwt(W_instr_L2_out_rsci_bdwt),
      .W_instr_L2_out_rsci_bcwt(W_instr_L2_out_rsci_bcwt),
      .W_instr_L2_out_rsci_ivld_run_sct(W_instr_L2_out_rsci_ivld_run_sct)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci_W_instr_L2_out_wait_dp
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci_W_instr_L2_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .W_instr_L2_out_rsci_oswt(W_instr_L2_out_rsci_oswt),
      .W_instr_L2_out_rsci_wen_comp(W_instr_L2_out_rsci_wen_comp),
      .W_instr_L2_out_rsci_biwt(W_instr_L2_out_rsci_biwt),
      .W_instr_L2_out_rsci_bdwt(W_instr_L2_out_rsci_bdwt),
      .W_instr_L2_out_rsci_bcwt(W_instr_L2_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci
    (
  clk, rst, W_instr_L1_out_rsc_dat, W_instr_L1_out_rsc_vld, W_instr_L1_out_rsc_rdy,
      run_wen, W_instr_L1_out_rsci_oswt, W_instr_L1_out_rsci_wen_comp, W_instr_L1_out_rsci_idat
);
  input clk;
  input rst;
  output [49:0] W_instr_L1_out_rsc_dat;
  output W_instr_L1_out_rsc_vld;
  input W_instr_L1_out_rsc_rdy;
  input run_wen;
  input W_instr_L1_out_rsci_oswt;
  output W_instr_L1_out_rsci_wen_comp;
  input [49:0] W_instr_L1_out_rsci_idat;


  // Interconnect Declarations
  wire W_instr_L1_out_rsci_irdy;
  wire W_instr_L1_out_rsci_biwt;
  wire W_instr_L1_out_rsci_bdwt;
  wire W_instr_L1_out_rsci_bcwt;
  wire W_instr_L1_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd33),
  .width(32'sd50)) W_instr_L1_out_rsci (
      .irdy(W_instr_L1_out_rsci_irdy),
      .ivld(W_instr_L1_out_rsci_ivld_run_sct),
      .idat(W_instr_L1_out_rsci_idat),
      .rdy(W_instr_L1_out_rsc_rdy),
      .vld(W_instr_L1_out_rsc_vld),
      .dat(W_instr_L1_out_rsc_dat)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci_W_instr_L1_out_wait_ctrl
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci_W_instr_L1_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .W_instr_L1_out_rsci_oswt(W_instr_L1_out_rsci_oswt),
      .W_instr_L1_out_rsci_irdy(W_instr_L1_out_rsci_irdy),
      .W_instr_L1_out_rsci_biwt(W_instr_L1_out_rsci_biwt),
      .W_instr_L1_out_rsci_bdwt(W_instr_L1_out_rsci_bdwt),
      .W_instr_L1_out_rsci_bcwt(W_instr_L1_out_rsci_bcwt),
      .W_instr_L1_out_rsci_ivld_run_sct(W_instr_L1_out_rsci_ivld_run_sct)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci_W_instr_L1_out_wait_dp
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci_W_instr_L1_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .W_instr_L1_out_rsci_oswt(W_instr_L1_out_rsci_oswt),
      .W_instr_L1_out_rsci_wen_comp(W_instr_L1_out_rsci_wen_comp),
      .W_instr_L1_out_rsci_biwt(W_instr_L1_out_rsci_biwt),
      .W_instr_L1_out_rsci_bdwt(W_instr_L1_out_rsci_bdwt),
      .W_instr_L1_out_rsci_bcwt(W_instr_L1_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci
    (
  clk, rst, I_instr_L3_out_rsc_dat, I_instr_L3_out_rsc_vld, I_instr_L3_out_rsc_rdy,
      run_wen, I_instr_L3_out_rsci_oswt, I_instr_L3_out_rsci_wen_comp, I_instr_L3_out_rsci_idat
);
  input clk;
  input rst;
  output [139:0] I_instr_L3_out_rsc_dat;
  output I_instr_L3_out_rsc_vld;
  input I_instr_L3_out_rsc_rdy;
  input run_wen;
  input I_instr_L3_out_rsci_oswt;
  output I_instr_L3_out_rsci_wen_comp;
  input [139:0] I_instr_L3_out_rsci_idat;


  // Interconnect Declarations
  wire I_instr_L3_out_rsci_irdy;
  wire I_instr_L3_out_rsci_biwt;
  wire I_instr_L3_out_rsci_bdwt;
  wire I_instr_L3_out_rsci_bcwt;
  wire I_instr_L3_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd32),
  .width(32'sd140)) I_instr_L3_out_rsci (
      .irdy(I_instr_L3_out_rsci_irdy),
      .ivld(I_instr_L3_out_rsci_ivld_run_sct),
      .idat(I_instr_L3_out_rsci_idat),
      .rdy(I_instr_L3_out_rsc_rdy),
      .vld(I_instr_L3_out_rsc_vld),
      .dat(I_instr_L3_out_rsc_dat)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci_I_instr_L3_out_wait_ctrl
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci_I_instr_L3_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .I_instr_L3_out_rsci_oswt(I_instr_L3_out_rsci_oswt),
      .I_instr_L3_out_rsci_irdy(I_instr_L3_out_rsci_irdy),
      .I_instr_L3_out_rsci_biwt(I_instr_L3_out_rsci_biwt),
      .I_instr_L3_out_rsci_bdwt(I_instr_L3_out_rsci_bdwt),
      .I_instr_L3_out_rsci_bcwt(I_instr_L3_out_rsci_bcwt),
      .I_instr_L3_out_rsci_ivld_run_sct(I_instr_L3_out_rsci_ivld_run_sct)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci_I_instr_L3_out_wait_dp
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci_I_instr_L3_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .I_instr_L3_out_rsci_oswt(I_instr_L3_out_rsci_oswt),
      .I_instr_L3_out_rsci_wen_comp(I_instr_L3_out_rsci_wen_comp),
      .I_instr_L3_out_rsci_biwt(I_instr_L3_out_rsci_biwt),
      .I_instr_L3_out_rsci_bdwt(I_instr_L3_out_rsci_bdwt),
      .I_instr_L3_out_rsci_bcwt(I_instr_L3_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci
    (
  clk, rst, I_instr_L2_out_rsc_dat, I_instr_L2_out_rsc_vld, I_instr_L2_out_rsc_rdy,
      run_wen, I_instr_L2_out_rsci_oswt, I_instr_L2_out_rsci_wen_comp, I_instr_L2_out_rsci_idat
);
  input clk;
  input rst;
  output [89:0] I_instr_L2_out_rsc_dat;
  output I_instr_L2_out_rsc_vld;
  input I_instr_L2_out_rsc_rdy;
  input run_wen;
  input I_instr_L2_out_rsci_oswt;
  output I_instr_L2_out_rsci_wen_comp;
  input [89:0] I_instr_L2_out_rsci_idat;


  // Interconnect Declarations
  wire I_instr_L2_out_rsci_irdy;
  wire I_instr_L2_out_rsci_biwt;
  wire I_instr_L2_out_rsci_bdwt;
  wire I_instr_L2_out_rsci_bcwt;
  wire I_instr_L2_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd31),
  .width(32'sd90)) I_instr_L2_out_rsci (
      .irdy(I_instr_L2_out_rsci_irdy),
      .ivld(I_instr_L2_out_rsci_ivld_run_sct),
      .idat(I_instr_L2_out_rsci_idat),
      .rdy(I_instr_L2_out_rsc_rdy),
      .vld(I_instr_L2_out_rsc_vld),
      .dat(I_instr_L2_out_rsc_dat)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci_I_instr_L2_out_wait_ctrl
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci_I_instr_L2_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .I_instr_L2_out_rsci_oswt(I_instr_L2_out_rsci_oswt),
      .I_instr_L2_out_rsci_irdy(I_instr_L2_out_rsci_irdy),
      .I_instr_L2_out_rsci_biwt(I_instr_L2_out_rsci_biwt),
      .I_instr_L2_out_rsci_bdwt(I_instr_L2_out_rsci_bdwt),
      .I_instr_L2_out_rsci_bcwt(I_instr_L2_out_rsci_bcwt),
      .I_instr_L2_out_rsci_ivld_run_sct(I_instr_L2_out_rsci_ivld_run_sct)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci_I_instr_L2_out_wait_dp
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci_I_instr_L2_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .I_instr_L2_out_rsci_oswt(I_instr_L2_out_rsci_oswt),
      .I_instr_L2_out_rsci_wen_comp(I_instr_L2_out_rsci_wen_comp),
      .I_instr_L2_out_rsci_biwt(I_instr_L2_out_rsci_biwt),
      .I_instr_L2_out_rsci_bdwt(I_instr_L2_out_rsci_bdwt),
      .I_instr_L2_out_rsci_bcwt(I_instr_L2_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci
    (
  clk, rst, I_instr_L1_out_rsc_dat, I_instr_L1_out_rsc_vld, I_instr_L1_out_rsc_rdy,
      run_wen, I_instr_L1_out_rsci_oswt, I_instr_L1_out_rsci_wen_comp, I_instr_L1_out_rsci_idat
);
  input clk;
  input rst;
  output [49:0] I_instr_L1_out_rsc_dat;
  output I_instr_L1_out_rsc_vld;
  input I_instr_L1_out_rsc_rdy;
  input run_wen;
  input I_instr_L1_out_rsci_oswt;
  output I_instr_L1_out_rsci_wen_comp;
  input [49:0] I_instr_L1_out_rsci_idat;


  // Interconnect Declarations
  wire I_instr_L1_out_rsci_irdy;
  wire I_instr_L1_out_rsci_biwt;
  wire I_instr_L1_out_rsci_bdwt;
  wire I_instr_L1_out_rsci_bcwt;
  wire I_instr_L1_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd30),
  .width(32'sd50)) I_instr_L1_out_rsci (
      .irdy(I_instr_L1_out_rsci_irdy),
      .ivld(I_instr_L1_out_rsci_ivld_run_sct),
      .idat(I_instr_L1_out_rsci_idat),
      .rdy(I_instr_L1_out_rsc_rdy),
      .vld(I_instr_L1_out_rsc_vld),
      .dat(I_instr_L1_out_rsc_dat)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci_I_instr_L1_out_wait_ctrl
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci_I_instr_L1_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .I_instr_L1_out_rsci_oswt(I_instr_L1_out_rsci_oswt),
      .I_instr_L1_out_rsci_irdy(I_instr_L1_out_rsci_irdy),
      .I_instr_L1_out_rsci_biwt(I_instr_L1_out_rsci_biwt),
      .I_instr_L1_out_rsci_bdwt(I_instr_L1_out_rsci_bdwt),
      .I_instr_L1_out_rsci_bcwt(I_instr_L1_out_rsci_bcwt),
      .I_instr_L1_out_rsci_ivld_run_sct(I_instr_L1_out_rsci_ivld_run_sct)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci_I_instr_L1_out_wait_dp
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci_I_instr_L1_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .I_instr_L1_out_rsci_oswt(I_instr_L1_out_rsci_oswt),
      .I_instr_L1_out_rsci_wen_comp(I_instr_L1_out_rsci_wen_comp),
      .I_instr_L1_out_rsci_biwt(I_instr_L1_out_rsci_biwt),
      .I_instr_L1_out_rsci_bdwt(I_instr_L1_out_rsci_bdwt),
      .I_instr_L1_out_rsci_bcwt(I_instr_L1_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci
    (
  clk, rst, O_instr_L3_out_rsc_dat, O_instr_L3_out_rsc_vld, O_instr_L3_out_rsc_rdy,
      run_wen, O_instr_L3_out_rsci_oswt, O_instr_L3_out_rsci_wen_comp, O_instr_L3_out_rsci_idat
);
  input clk;
  input rst;
  output [139:0] O_instr_L3_out_rsc_dat;
  output O_instr_L3_out_rsc_vld;
  input O_instr_L3_out_rsc_rdy;
  input run_wen;
  input O_instr_L3_out_rsci_oswt;
  output O_instr_L3_out_rsci_wen_comp;
  input [139:0] O_instr_L3_out_rsci_idat;


  // Interconnect Declarations
  wire O_instr_L3_out_rsci_irdy;
  wire O_instr_L3_out_rsci_biwt;
  wire O_instr_L3_out_rsci_bdwt;
  wire O_instr_L3_out_rsci_bcwt;
  wire O_instr_L3_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd29),
  .width(32'sd140)) O_instr_L3_out_rsci (
      .irdy(O_instr_L3_out_rsci_irdy),
      .ivld(O_instr_L3_out_rsci_ivld_run_sct),
      .idat(O_instr_L3_out_rsci_idat),
      .rdy(O_instr_L3_out_rsc_rdy),
      .vld(O_instr_L3_out_rsc_vld),
      .dat(O_instr_L3_out_rsc_dat)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci_O_instr_L3_out_wait_ctrl
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci_O_instr_L3_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .O_instr_L3_out_rsci_oswt(O_instr_L3_out_rsci_oswt),
      .O_instr_L3_out_rsci_irdy(O_instr_L3_out_rsci_irdy),
      .O_instr_L3_out_rsci_biwt(O_instr_L3_out_rsci_biwt),
      .O_instr_L3_out_rsci_bdwt(O_instr_L3_out_rsci_bdwt),
      .O_instr_L3_out_rsci_bcwt(O_instr_L3_out_rsci_bcwt),
      .O_instr_L3_out_rsci_ivld_run_sct(O_instr_L3_out_rsci_ivld_run_sct)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci_O_instr_L3_out_wait_dp
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci_O_instr_L3_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .O_instr_L3_out_rsci_oswt(O_instr_L3_out_rsci_oswt),
      .O_instr_L3_out_rsci_wen_comp(O_instr_L3_out_rsci_wen_comp),
      .O_instr_L3_out_rsci_biwt(O_instr_L3_out_rsci_biwt),
      .O_instr_L3_out_rsci_bdwt(O_instr_L3_out_rsci_bdwt),
      .O_instr_L3_out_rsci_bcwt(O_instr_L3_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci
    (
  clk, rst, O_instr_L2_out_rsc_dat, O_instr_L2_out_rsc_vld, O_instr_L2_out_rsc_rdy,
      run_wen, O_instr_L2_out_rsci_oswt, O_instr_L2_out_rsci_wen_comp, O_instr_L2_out_rsci_idat
);
  input clk;
  input rst;
  output [89:0] O_instr_L2_out_rsc_dat;
  output O_instr_L2_out_rsc_vld;
  input O_instr_L2_out_rsc_rdy;
  input run_wen;
  input O_instr_L2_out_rsci_oswt;
  output O_instr_L2_out_rsci_wen_comp;
  input [89:0] O_instr_L2_out_rsci_idat;


  // Interconnect Declarations
  wire O_instr_L2_out_rsci_irdy;
  wire O_instr_L2_out_rsci_biwt;
  wire O_instr_L2_out_rsci_bdwt;
  wire O_instr_L2_out_rsci_bcwt;
  wire O_instr_L2_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd28),
  .width(32'sd90)) O_instr_L2_out_rsci (
      .irdy(O_instr_L2_out_rsci_irdy),
      .ivld(O_instr_L2_out_rsci_ivld_run_sct),
      .idat(O_instr_L2_out_rsci_idat),
      .rdy(O_instr_L2_out_rsc_rdy),
      .vld(O_instr_L2_out_rsc_vld),
      .dat(O_instr_L2_out_rsc_dat)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci_O_instr_L2_out_wait_ctrl
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci_O_instr_L2_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .O_instr_L2_out_rsci_oswt(O_instr_L2_out_rsci_oswt),
      .O_instr_L2_out_rsci_irdy(O_instr_L2_out_rsci_irdy),
      .O_instr_L2_out_rsci_biwt(O_instr_L2_out_rsci_biwt),
      .O_instr_L2_out_rsci_bdwt(O_instr_L2_out_rsci_bdwt),
      .O_instr_L2_out_rsci_bcwt(O_instr_L2_out_rsci_bcwt),
      .O_instr_L2_out_rsci_ivld_run_sct(O_instr_L2_out_rsci_ivld_run_sct)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci_O_instr_L2_out_wait_dp
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci_O_instr_L2_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .O_instr_L2_out_rsci_oswt(O_instr_L2_out_rsci_oswt),
      .O_instr_L2_out_rsci_wen_comp(O_instr_L2_out_rsci_wen_comp),
      .O_instr_L2_out_rsci_biwt(O_instr_L2_out_rsci_biwt),
      .O_instr_L2_out_rsci_bdwt(O_instr_L2_out_rsci_bdwt),
      .O_instr_L2_out_rsci_bcwt(O_instr_L2_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci
    (
  clk, rst, O_instr_L1_out_rsc_dat, O_instr_L1_out_rsc_vld, O_instr_L1_out_rsc_rdy,
      run_wen, O_instr_L1_out_rsci_oswt, O_instr_L1_out_rsci_wen_comp, O_instr_L1_out_rsci_idat
);
  input clk;
  input rst;
  output [49:0] O_instr_L1_out_rsc_dat;
  output O_instr_L1_out_rsc_vld;
  input O_instr_L1_out_rsc_rdy;
  input run_wen;
  input O_instr_L1_out_rsci_oswt;
  output O_instr_L1_out_rsci_wen_comp;
  input [49:0] O_instr_L1_out_rsci_idat;


  // Interconnect Declarations
  wire O_instr_L1_out_rsci_irdy;
  wire O_instr_L1_out_rsci_biwt;
  wire O_instr_L1_out_rsci_bdwt;
  wire O_instr_L1_out_rsci_bcwt;
  wire O_instr_L1_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd27),
  .width(32'sd50)) O_instr_L1_out_rsci (
      .irdy(O_instr_L1_out_rsci_irdy),
      .ivld(O_instr_L1_out_rsci_ivld_run_sct),
      .idat(O_instr_L1_out_rsci_idat),
      .rdy(O_instr_L1_out_rsc_rdy),
      .vld(O_instr_L1_out_rsc_vld),
      .dat(O_instr_L1_out_rsc_dat)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci_O_instr_L1_out_wait_ctrl
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci_O_instr_L1_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .O_instr_L1_out_rsci_oswt(O_instr_L1_out_rsci_oswt),
      .O_instr_L1_out_rsci_irdy(O_instr_L1_out_rsci_irdy),
      .O_instr_L1_out_rsci_biwt(O_instr_L1_out_rsci_biwt),
      .O_instr_L1_out_rsci_bdwt(O_instr_L1_out_rsci_bdwt),
      .O_instr_L1_out_rsci_bcwt(O_instr_L1_out_rsci_bcwt),
      .O_instr_L1_out_rsci_ivld_run_sct(O_instr_L1_out_rsci_ivld_run_sct)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci_O_instr_L1_out_wait_dp
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci_O_instr_L1_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .O_instr_L1_out_rsci_oswt(O_instr_L1_out_rsci_oswt),
      .O_instr_L1_out_rsci_wen_comp(O_instr_L1_out_rsci_wen_comp),
      .O_instr_L1_out_rsci_biwt(O_instr_L1_out_rsci_biwt),
      .O_instr_L1_out_rsci_bdwt(O_instr_L1_out_rsci_bdwt),
      .O_instr_L1_out_rsci_bcwt(O_instr_L1_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_layer_instruction_in_rsci
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_layer_instruction_in_rsci
    (
  clk, rst, layer_instruction_in_rsc_dat, layer_instruction_in_rsc_vld, layer_instruction_in_rsc_rdy,
      run_wen, layer_instruction_in_rsci_oswt, layer_instruction_in_rsci_wen_comp,
      layer_instruction_in_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [484:0] layer_instruction_in_rsc_dat;
  input layer_instruction_in_rsc_vld;
  output layer_instruction_in_rsc_rdy;
  input run_wen;
  input layer_instruction_in_rsci_oswt;
  output layer_instruction_in_rsci_wen_comp;
  output [484:0] layer_instruction_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire layer_instruction_in_rsci_biwt;
  wire layer_instruction_in_rsci_bdwt;
  wire layer_instruction_in_rsci_bcwt;
  wire layer_instruction_in_rsci_irdy_run_sct;
  wire layer_instruction_in_rsci_ivld;
  wire [484:0] layer_instruction_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd26),
  .width(32'sd485)) layer_instruction_in_rsci (
      .rdy(layer_instruction_in_rsc_rdy),
      .vld(layer_instruction_in_rsc_vld),
      .dat(layer_instruction_in_rsc_dat),
      .irdy(layer_instruction_in_rsci_irdy_run_sct),
      .ivld(layer_instruction_in_rsci_ivld),
      .idat(layer_instruction_in_rsci_idat)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_layer_instruction_in_rsci_layer_instruction_in_wait_ctrl
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_layer_instruction_in_rsci_layer_instruction_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .layer_instruction_in_rsci_oswt(layer_instruction_in_rsci_oswt),
      .layer_instruction_in_rsci_biwt(layer_instruction_in_rsci_biwt),
      .layer_instruction_in_rsci_bdwt(layer_instruction_in_rsci_bdwt),
      .layer_instruction_in_rsci_bcwt(layer_instruction_in_rsci_bcwt),
      .layer_instruction_in_rsci_irdy_run_sct(layer_instruction_in_rsci_irdy_run_sct),
      .layer_instruction_in_rsci_ivld(layer_instruction_in_rsci_ivld)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_layer_instruction_in_rsci_layer_instruction_in_wait_dp
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_layer_instruction_in_rsci_layer_instruction_in_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .layer_instruction_in_rsci_oswt(layer_instruction_in_rsci_oswt),
      .layer_instruction_in_rsci_wen_comp(layer_instruction_in_rsci_wen_comp),
      .layer_instruction_in_rsci_idat_mxwt(layer_instruction_in_rsci_idat_mxwt),
      .layer_instruction_in_rsci_biwt(layer_instruction_in_rsci_biwt),
      .layer_instruction_in_rsci_bdwt(layer_instruction_in_rsci_bdwt),
      .layer_instruction_in_rsci_bcwt(layer_instruction_in_rsci_bcwt),
      .layer_instruction_in_rsci_idat(layer_instruction_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_instr_in_rsci
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_instr_in_rsci
    (
  clk, rst, W_instr_in_rsc_dat, W_instr_in_rsc_vld, W_instr_in_rsc_rdy, run_wen,
      W_instr_in_rsci_oswt, W_instr_in_rsci_wen_comp, W_instr_in_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [49:0] W_instr_in_rsc_dat;
  input W_instr_in_rsc_vld;
  output W_instr_in_rsc_rdy;
  input run_wen;
  input W_instr_in_rsci_oswt;
  output W_instr_in_rsci_wen_comp;
  output [49:0] W_instr_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire W_instr_in_rsci_biwt;
  wire W_instr_in_rsci_bdwt;
  wire W_instr_in_rsci_bcwt;
  wire W_instr_in_rsci_irdy_run_sct;
  wire W_instr_in_rsci_ivld;
  wire [49:0] W_instr_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd75),
  .width(32'sd50)) W_instr_in_rsci (
      .rdy(W_instr_in_rsc_rdy),
      .vld(W_instr_in_rsc_vld),
      .dat(W_instr_in_rsc_dat),
      .irdy(W_instr_in_rsci_irdy_run_sct),
      .ivld(W_instr_in_rsci_ivld),
      .idat(W_instr_in_rsci_idat)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_instr_in_rsci_W_instr_in_wait_ctrl
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_instr_in_rsci_W_instr_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .W_instr_in_rsci_oswt(W_instr_in_rsci_oswt),
      .W_instr_in_rsci_biwt(W_instr_in_rsci_biwt),
      .W_instr_in_rsci_bdwt(W_instr_in_rsci_bdwt),
      .W_instr_in_rsci_bcwt(W_instr_in_rsci_bcwt),
      .W_instr_in_rsci_irdy_run_sct(W_instr_in_rsci_irdy_run_sct),
      .W_instr_in_rsci_ivld(W_instr_in_rsci_ivld)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_instr_in_rsci_W_instr_in_wait_dp
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_instr_in_rsci_W_instr_in_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .W_instr_in_rsci_oswt(W_instr_in_rsci_oswt),
      .W_instr_in_rsci_wen_comp(W_instr_in_rsci_wen_comp),
      .W_instr_in_rsci_idat_mxwt(W_instr_in_rsci_idat_mxwt),
      .W_instr_in_rsci_biwt(W_instr_in_rsci_biwt),
      .W_instr_in_rsci_bdwt(W_instr_in_rsci_bdwt),
      .W_instr_in_rsci_bcwt(W_instr_in_rsci_bcwt),
      .W_instr_in_rsci_idat(W_instr_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_instr_in_rsci
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_instr_in_rsci
    (
  clk, rst, I_instr_in_rsc_dat, I_instr_in_rsc_vld, I_instr_in_rsc_rdy, run_wen,
      I_instr_in_rsci_oswt, I_instr_in_rsci_wen_comp, I_instr_in_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [49:0] I_instr_in_rsc_dat;
  input I_instr_in_rsc_vld;
  output I_instr_in_rsc_rdy;
  input run_wen;
  input I_instr_in_rsci_oswt;
  output I_instr_in_rsci_wen_comp;
  output [49:0] I_instr_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire I_instr_in_rsci_biwt;
  wire I_instr_in_rsci_bdwt;
  wire I_instr_in_rsci_bcwt;
  wire I_instr_in_rsci_irdy_run_sct;
  wire I_instr_in_rsci_ivld;
  wire [49:0] I_instr_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd74),
  .width(32'sd50)) I_instr_in_rsci (
      .rdy(I_instr_in_rsc_rdy),
      .vld(I_instr_in_rsc_vld),
      .dat(I_instr_in_rsc_dat),
      .irdy(I_instr_in_rsci_irdy_run_sct),
      .ivld(I_instr_in_rsci_ivld),
      .idat(I_instr_in_rsci_idat)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_instr_in_rsci_I_instr_in_wait_ctrl
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_instr_in_rsci_I_instr_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .I_instr_in_rsci_oswt(I_instr_in_rsci_oswt),
      .I_instr_in_rsci_biwt(I_instr_in_rsci_biwt),
      .I_instr_in_rsci_bdwt(I_instr_in_rsci_bdwt),
      .I_instr_in_rsci_bcwt(I_instr_in_rsci_bcwt),
      .I_instr_in_rsci_irdy_run_sct(I_instr_in_rsci_irdy_run_sct),
      .I_instr_in_rsci_ivld(I_instr_in_rsci_ivld)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_instr_in_rsci_I_instr_in_wait_dp
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_instr_in_rsci_I_instr_in_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .I_instr_in_rsci_oswt(I_instr_in_rsci_oswt),
      .I_instr_in_rsci_wen_comp(I_instr_in_rsci_wen_comp),
      .I_instr_in_rsci_idat_mxwt(I_instr_in_rsci_idat_mxwt),
      .I_instr_in_rsci_biwt(I_instr_in_rsci_biwt),
      .I_instr_in_rsci_bdwt(I_instr_in_rsci_bdwt),
      .I_instr_in_rsci_bcwt(I_instr_in_rsci_bcwt),
      .I_instr_in_rsci_idat(I_instr_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_instr_in_rsci
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_instr_in_rsci
    (
  clk, rst, O_instr_in_rsc_dat, O_instr_in_rsc_vld, O_instr_in_rsc_rdy, run_wen,
      O_instr_in_rsci_oswt, O_instr_in_rsci_wen_comp, O_instr_in_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [49:0] O_instr_in_rsc_dat;
  input O_instr_in_rsc_vld;
  output O_instr_in_rsc_rdy;
  input run_wen;
  input O_instr_in_rsci_oswt;
  output O_instr_in_rsci_wen_comp;
  output [49:0] O_instr_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire O_instr_in_rsci_biwt;
  wire O_instr_in_rsci_bdwt;
  wire O_instr_in_rsci_bcwt;
  wire O_instr_in_rsci_irdy_run_sct;
  wire O_instr_in_rsci_ivld;
  wire [49:0] O_instr_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd73),
  .width(32'sd50)) O_instr_in_rsci (
      .rdy(O_instr_in_rsc_rdy),
      .vld(O_instr_in_rsc_vld),
      .dat(O_instr_in_rsc_dat),
      .irdy(O_instr_in_rsci_irdy_run_sct),
      .ivld(O_instr_in_rsci_ivld),
      .idat(O_instr_in_rsci_idat)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_instr_in_rsci_O_instr_in_wait_ctrl
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_instr_in_rsci_O_instr_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .O_instr_in_rsci_oswt(O_instr_in_rsci_oswt),
      .O_instr_in_rsci_biwt(O_instr_in_rsci_biwt),
      .O_instr_in_rsci_bdwt(O_instr_in_rsci_bdwt),
      .O_instr_in_rsci_bcwt(O_instr_in_rsci_bcwt),
      .O_instr_in_rsci_irdy_run_sct(O_instr_in_rsci_irdy_run_sct),
      .O_instr_in_rsci_ivld(O_instr_in_rsci_ivld)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_instr_in_rsci_O_instr_in_wait_dp
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_instr_in_rsci_O_instr_in_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .O_instr_in_rsci_oswt(O_instr_in_rsci_oswt),
      .O_instr_in_rsci_wen_comp(O_instr_in_rsci_wen_comp),
      .O_instr_in_rsci_idat_mxwt(O_instr_in_rsci_idat_mxwt),
      .O_instr_in_rsci_biwt(O_instr_in_rsci_biwt),
      .O_instr_in_rsci_bdwt(O_instr_in_rsci_bdwt),
      .O_instr_in_rsci_bcwt(O_instr_in_rsci_bcwt),
      .O_instr_in_rsci_idat(O_instr_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_wr_data_zero_guard_rsci
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_wr_data_zero_guard_rsci
    (
  clk, rst, wr_data_zero_guard_rsc_dat, wr_data_zero_guard_rsc_vld, wr_data_zero_guard_rsc_rdy,
      run_wen, run_wten, wr_data_zero_guard_rsci_oswt, wr_data_zero_guard_rsci_ivld_mxwt,
      wr_data_zero_guard_rsci_idat_mxwt
);
  input clk;
  input rst;
  input wr_data_zero_guard_rsc_dat;
  input wr_data_zero_guard_rsc_vld;
  output wr_data_zero_guard_rsc_rdy;
  input run_wen;
  input run_wten;
  input wr_data_zero_guard_rsci_oswt;
  output wr_data_zero_guard_rsci_ivld_mxwt;
  output wr_data_zero_guard_rsci_idat_mxwt;


  // Interconnect Declarations
  wire wr_data_zero_guard_rsci_biwt;
  wire wr_data_zero_guard_rsci_bdwt;
  wire wr_data_zero_guard_rsci_ivld;
  wire wr_data_zero_guard_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd72),
  .width(32'sd1)) wr_data_zero_guard_rsci (
      .rdy(wr_data_zero_guard_rsc_rdy),
      .vld(wr_data_zero_guard_rsc_vld),
      .dat(wr_data_zero_guard_rsc_dat),
      .irdy(wr_data_zero_guard_rsci_biwt),
      .ivld(wr_data_zero_guard_rsci_ivld),
      .idat(wr_data_zero_guard_rsci_idat)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_wr_data_zero_guard_rsci_wr_data_zero_guard_wait_ctrl
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_wr_data_zero_guard_rsci_wr_data_zero_guard_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .wr_data_zero_guard_rsci_oswt(wr_data_zero_guard_rsci_oswt),
      .wr_data_zero_guard_rsci_biwt(wr_data_zero_guard_rsci_biwt),
      .wr_data_zero_guard_rsci_bdwt(wr_data_zero_guard_rsci_bdwt)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_wr_data_zero_guard_rsci_wr_data_zero_guard_wait_dp
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_wr_data_zero_guard_rsci_wr_data_zero_guard_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .wr_data_zero_guard_rsci_ivld_mxwt(wr_data_zero_guard_rsci_ivld_mxwt),
      .wr_data_zero_guard_rsci_idat_mxwt(wr_data_zero_guard_rsci_idat_mxwt),
      .wr_data_zero_guard_rsci_biwt(wr_data_zero_guard_rsci_biwt),
      .wr_data_zero_guard_rsci_bdwt(wr_data_zero_guard_rsci_bdwt),
      .wr_data_zero_guard_rsci_ivld(wr_data_zero_guard_rsci_ivld),
      .wr_data_zero_guard_rsci_idat(wr_data_zero_guard_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_wr_data_rsci
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_wr_data_rsci
    (
  clk, rst, W_wr_data_rsc_dat, W_wr_data_rsc_vld, W_wr_data_rsc_rdy, run_wen, run_wten,
      W_wr_data_rsci_oswt, W_wr_data_rsci_ivld_mxwt, W_wr_data_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [15:0] W_wr_data_rsc_dat;
  input W_wr_data_rsc_vld;
  output W_wr_data_rsc_rdy;
  input run_wen;
  input run_wten;
  input W_wr_data_rsci_oswt;
  output W_wr_data_rsci_ivld_mxwt;
  output [15:0] W_wr_data_rsci_idat_mxwt;


  // Interconnect Declarations
  wire W_wr_data_rsci_biwt;
  wire W_wr_data_rsci_bdwt;
  wire W_wr_data_rsci_ivld;
  wire [15:0] W_wr_data_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd71),
  .width(32'sd16)) W_wr_data_rsci (
      .rdy(W_wr_data_rsc_rdy),
      .vld(W_wr_data_rsc_vld),
      .dat(W_wr_data_rsc_dat),
      .irdy(W_wr_data_rsci_biwt),
      .ivld(W_wr_data_rsci_ivld),
      .idat(W_wr_data_rsci_idat)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_wr_data_rsci_W_wr_data_wait_ctrl
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_wr_data_rsci_W_wr_data_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .W_wr_data_rsci_oswt(W_wr_data_rsci_oswt),
      .W_wr_data_rsci_biwt(W_wr_data_rsci_biwt),
      .W_wr_data_rsci_bdwt(W_wr_data_rsci_bdwt)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_wr_data_rsci_W_wr_data_wait_dp
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_wr_data_rsci_W_wr_data_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .W_wr_data_rsci_ivld_mxwt(W_wr_data_rsci_ivld_mxwt),
      .W_wr_data_rsci_idat_mxwt(W_wr_data_rsci_idat_mxwt),
      .W_wr_data_rsci_biwt(W_wr_data_rsci_biwt),
      .W_wr_data_rsci_bdwt(W_wr_data_rsci_bdwt),
      .W_wr_data_rsci_ivld(W_wr_data_rsci_ivld),
      .W_wr_data_rsci_idat(W_wr_data_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_wr_data_rsci
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_wr_data_rsci
    (
  clk, rst, I_wr_data_rsc_dat, I_wr_data_rsc_vld, I_wr_data_rsc_rdy, run_wen, run_wten,
      I_wr_data_rsci_oswt, I_wr_data_rsci_ivld_mxwt, I_wr_data_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [15:0] I_wr_data_rsc_dat;
  input I_wr_data_rsc_vld;
  output I_wr_data_rsc_rdy;
  input run_wen;
  input run_wten;
  input I_wr_data_rsci_oswt;
  output I_wr_data_rsci_ivld_mxwt;
  output [15:0] I_wr_data_rsci_idat_mxwt;


  // Interconnect Declarations
  wire I_wr_data_rsci_biwt;
  wire I_wr_data_rsci_bdwt;
  wire I_wr_data_rsci_ivld;
  wire [15:0] I_wr_data_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd70),
  .width(32'sd16)) I_wr_data_rsci (
      .rdy(I_wr_data_rsc_rdy),
      .vld(I_wr_data_rsc_vld),
      .dat(I_wr_data_rsc_dat),
      .irdy(I_wr_data_rsci_biwt),
      .ivld(I_wr_data_rsci_ivld),
      .idat(I_wr_data_rsci_idat)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_wr_data_rsci_I_wr_data_wait_ctrl
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_wr_data_rsci_I_wr_data_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .I_wr_data_rsci_oswt(I_wr_data_rsci_oswt),
      .I_wr_data_rsci_biwt(I_wr_data_rsci_biwt),
      .I_wr_data_rsci_bdwt(I_wr_data_rsci_bdwt)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_wr_data_rsci_I_wr_data_wait_dp
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_wr_data_rsci_I_wr_data_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .I_wr_data_rsci_ivld_mxwt(I_wr_data_rsci_ivld_mxwt),
      .I_wr_data_rsci_idat_mxwt(I_wr_data_rsci_idat_mxwt),
      .I_wr_data_rsci_biwt(I_wr_data_rsci_biwt),
      .I_wr_data_rsci_bdwt(I_wr_data_rsci_bdwt),
      .I_wr_data_rsci_ivld(I_wr_data_rsci_ivld),
      .I_wr_data_rsci_idat(I_wr_data_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_rd_data_rsci
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_rd_data_rsci
    (
  clk, rst, O_rd_data_rsc_dat, O_rd_data_rsc_vld, O_rd_data_rsc_rdy, run_wen, run_wten,
      O_rd_data_rsci_oswt, O_rd_data_rsci_irdy_mxwt, O_rd_data_rsci_idat
);
  input clk;
  input rst;
  output [15:0] O_rd_data_rsc_dat;
  output O_rd_data_rsc_vld;
  input O_rd_data_rsc_rdy;
  input run_wen;
  input run_wten;
  input O_rd_data_rsci_oswt;
  output O_rd_data_rsci_irdy_mxwt;
  input [15:0] O_rd_data_rsci_idat;


  // Interconnect Declarations
  wire O_rd_data_rsci_irdy;
  wire O_rd_data_rsci_biwt;
  wire O_rd_data_rsci_bdwt;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd69),
  .width(32'sd16)) O_rd_data_rsci (
      .irdy(O_rd_data_rsci_irdy),
      .ivld(O_rd_data_rsci_biwt),
      .idat(O_rd_data_rsci_idat),
      .rdy(O_rd_data_rsc_rdy),
      .vld(O_rd_data_rsc_vld),
      .dat(O_rd_data_rsc_dat)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_rd_data_rsci_O_rd_data_wait_ctrl
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_rd_data_rsci_O_rd_data_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .O_rd_data_rsci_oswt(O_rd_data_rsci_oswt),
      .O_rd_data_rsci_biwt(O_rd_data_rsci_biwt),
      .O_rd_data_rsci_bdwt(O_rd_data_rsci_bdwt)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_rd_data_rsci_O_rd_data_wait_dp
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_rd_data_rsci_O_rd_data_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .O_rd_data_rsci_irdy_mxwt(O_rd_data_rsci_irdy_mxwt),
      .O_rd_data_rsci_irdy(O_rd_data_rsci_irdy),
      .O_rd_data_rsci_biwt(O_rd_data_rsci_biwt),
      .O_rd_data_rsci_bdwt(O_rd_data_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_wr_data_rsci
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_wr_data_rsci
    (
  clk, rst, O_wr_data_rsc_dat, O_wr_data_rsc_vld, O_wr_data_rsc_rdy, run_wen, O_wr_data_rsci_oswt,
      run_wten, O_wr_data_rsci_ivld_mxwt, O_wr_data_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [15:0] O_wr_data_rsc_dat;
  input O_wr_data_rsc_vld;
  output O_wr_data_rsc_rdy;
  input run_wen;
  input O_wr_data_rsci_oswt;
  input run_wten;
  output O_wr_data_rsci_ivld_mxwt;
  output [15:0] O_wr_data_rsci_idat_mxwt;


  // Interconnect Declarations
  wire O_wr_data_rsci_biwt;
  wire O_wr_data_rsci_bdwt;
  wire O_wr_data_rsci_ivld;
  wire [15:0] O_wr_data_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd68),
  .width(32'sd16)) O_wr_data_rsci (
      .rdy(O_wr_data_rsc_rdy),
      .vld(O_wr_data_rsc_vld),
      .dat(O_wr_data_rsc_dat),
      .irdy(O_wr_data_rsci_biwt),
      .ivld(O_wr_data_rsci_ivld),
      .idat(O_wr_data_rsci_idat)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_wr_data_rsci_O_wr_data_wait_ctrl
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_wr_data_rsci_O_wr_data_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .O_wr_data_rsci_oswt(O_wr_data_rsci_oswt),
      .run_wten(run_wten),
      .O_wr_data_rsci_biwt(O_wr_data_rsci_biwt),
      .O_wr_data_rsci_bdwt(O_wr_data_rsci_bdwt)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_wr_data_rsci_O_wr_data_wait_dp
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_wr_data_rsci_O_wr_data_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .O_wr_data_rsci_ivld_mxwt(O_wr_data_rsci_ivld_mxwt),
      .O_wr_data_rsci_idat_mxwt(O_wr_data_rsci_idat_mxwt),
      .O_wr_data_rsci_biwt(O_wr_data_rsci_biwt),
      .O_wr_data_rsci_bdwt(O_wr_data_rsci_bdwt),
      .O_wr_data_rsci_ivld(O_wr_data_rsci_ivld),
      .O_wr_data_rsci_idat(O_wr_data_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run
    (
  clk, rst, layer_instruction_in_rsc_dat, layer_instruction_in_rsc_vld, layer_instruction_in_rsc_rdy,
      O_instr_L1_out_rsc_dat, O_instr_L1_out_rsc_vld, O_instr_L1_out_rsc_rdy, O_instr_L2_out_rsc_dat,
      O_instr_L2_out_rsc_vld, O_instr_L2_out_rsc_rdy, O_instr_L3_out_rsc_dat, O_instr_L3_out_rsc_vld,
      O_instr_L3_out_rsc_rdy, I_instr_L1_out_rsc_dat, I_instr_L1_out_rsc_vld, I_instr_L1_out_rsc_rdy,
      I_instr_L2_out_rsc_dat, I_instr_L2_out_rsc_vld, I_instr_L2_out_rsc_rdy, I_instr_L3_out_rsc_dat,
      I_instr_L3_out_rsc_vld, I_instr_L3_out_rsc_rdy, W_instr_L1_out_rsc_dat, W_instr_L1_out_rsc_vld,
      W_instr_L1_out_rsc_rdy, W_instr_L2_out_rsc_dat, W_instr_L2_out_rsc_vld, W_instr_L2_out_rsc_rdy,
      W_instr_L3_out_rsc_dat, W_instr_L3_out_rsc_vld, W_instr_L3_out_rsc_rdy, W_tiling_unit_L3_run_cmp_loops_bound_rsc_dat,
      W_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat, W_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat,
      W_tiling_unit_L3_run_cmp_instr_bound_rsc_z, W_tiling_unit_L3_run_cmp_instr_tile_rsc_z,
      W_tiling_unit_L3_run_cmp_ccs_ccore_start_rsc_dat, W_tiling_unit_L3_run_cmp_ccs_ccore_en,
      ensig_cgo_iro_1, CGHpart_irsig_1, W_tiling_unit_L2_run_cmp_loops_bound_rsc_dat,
      W_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat, W_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat,
      W_tiling_unit_L2_run_cmp_tile_size_out_rsc_z, W_tiling_unit_L2_run_cmp_instr_bound_rsc_z,
      W_tiling_unit_L2_run_cmp_instr_tile_rsc_z, W_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat,
      W_tiling_unit_L2_run_cmp_ccs_ccore_en, O_tiling_unit_L3_run_cmp_loops_bound_rsc_dat,
      O_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat, O_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat,
      O_tiling_unit_L3_run_cmp_instr_bound_rsc_z, O_tiling_unit_L3_run_cmp_instr_tile_rsc_z,
      O_tiling_unit_L3_run_cmp_ccs_ccore_en, O_tiling_unit_L2_run_cmp_loops_bound_rsc_dat,
      O_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat, O_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat,
      O_tiling_unit_L2_run_cmp_tile_size_out_rsc_z, O_tiling_unit_L2_run_cmp_instr_bound_rsc_z,
      O_tiling_unit_L2_run_cmp_instr_tile_rsc_z, O_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat,
      O_tiling_unit_L2_run_cmp_ccs_ccore_en, O_tiling_unit_L1_run_cmp_loops_bound_rsc_dat,
      O_tiling_unit_L1_run_cmp_loops_relevancy_rsc_dat, O_tiling_unit_L1_run_cmp_tile_size_in_rsc_dat,
      O_tiling_unit_L1_run_cmp_tile_size_out_rsc_z, O_tiling_unit_L1_run_cmp_instr_bound_rsc_z,
      O_tiling_unit_L1_run_cmp_instr_tile_rsc_z, O_tiling_unit_L1_run_cmp_ccs_ccore_start_rsc_dat,
      O_tiling_unit_L1_run_cmp_ccs_ccore_en
);
  input clk;
  input rst;
  input [484:0] layer_instruction_in_rsc_dat;
  input layer_instruction_in_rsc_vld;
  output layer_instruction_in_rsc_rdy;
  output [49:0] O_instr_L1_out_rsc_dat;
  output O_instr_L1_out_rsc_vld;
  input O_instr_L1_out_rsc_rdy;
  output [89:0] O_instr_L2_out_rsc_dat;
  output O_instr_L2_out_rsc_vld;
  input O_instr_L2_out_rsc_rdy;
  output [139:0] O_instr_L3_out_rsc_dat;
  output O_instr_L3_out_rsc_vld;
  input O_instr_L3_out_rsc_rdy;
  output [49:0] I_instr_L1_out_rsc_dat;
  output I_instr_L1_out_rsc_vld;
  input I_instr_L1_out_rsc_rdy;
  output [89:0] I_instr_L2_out_rsc_dat;
  output I_instr_L2_out_rsc_vld;
  input I_instr_L2_out_rsc_rdy;
  output [139:0] I_instr_L3_out_rsc_dat;
  output I_instr_L3_out_rsc_vld;
  input I_instr_L3_out_rsc_rdy;
  output [49:0] W_instr_L1_out_rsc_dat;
  output W_instr_L1_out_rsc_vld;
  input W_instr_L1_out_rsc_rdy;
  output [109:0] W_instr_L2_out_rsc_dat;
  output W_instr_L2_out_rsc_vld;
  input W_instr_L2_out_rsc_rdy;
  output [159:0] W_instr_L3_out_rsc_dat;
  output W_instr_L3_out_rsc_vld;
  input W_instr_L3_out_rsc_rdy;
  output [79:0] W_tiling_unit_L3_run_cmp_loops_bound_rsc_dat;
  output [4:0] W_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat;
  output [15:0] W_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat;
  input [79:0] W_tiling_unit_L3_run_cmp_instr_bound_rsc_z;
  input [79:0] W_tiling_unit_L3_run_cmp_instr_tile_rsc_z;
  output W_tiling_unit_L3_run_cmp_ccs_ccore_start_rsc_dat;
  output W_tiling_unit_L3_run_cmp_ccs_ccore_en;
  input ensig_cgo_iro_1;
  output CGHpart_irsig_1;
  output [54:0] W_tiling_unit_L2_run_cmp_loops_bound_rsc_dat;
  output [4:0] W_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat;
  output [10:0] W_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat;
  input [10:0] W_tiling_unit_L2_run_cmp_tile_size_out_rsc_z;
  input [54:0] W_tiling_unit_L2_run_cmp_instr_bound_rsc_z;
  input [54:0] W_tiling_unit_L2_run_cmp_instr_tile_rsc_z;
  output W_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat;
  output W_tiling_unit_L2_run_cmp_ccs_ccore_en;
  output [69:0] O_tiling_unit_L3_run_cmp_loops_bound_rsc_dat;
  output [4:0] O_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat;
  output [13:0] O_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat;
  input [69:0] O_tiling_unit_L3_run_cmp_instr_bound_rsc_z;
  input [69:0] O_tiling_unit_L3_run_cmp_instr_tile_rsc_z;
  output O_tiling_unit_L3_run_cmp_ccs_ccore_en;
  output [44:0] O_tiling_unit_L2_run_cmp_loops_bound_rsc_dat;
  output [4:0] O_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat;
  output [8:0] O_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat;
  input [8:0] O_tiling_unit_L2_run_cmp_tile_size_out_rsc_z;
  input [44:0] O_tiling_unit_L2_run_cmp_instr_bound_rsc_z;
  input [44:0] O_tiling_unit_L2_run_cmp_instr_tile_rsc_z;
  output O_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat;
  output O_tiling_unit_L2_run_cmp_ccs_ccore_en;
  output [24:0] O_tiling_unit_L1_run_cmp_loops_bound_rsc_dat;
  output [4:0] O_tiling_unit_L1_run_cmp_loops_relevancy_rsc_dat;
  output [4:0] O_tiling_unit_L1_run_cmp_tile_size_in_rsc_dat;
  input [4:0] O_tiling_unit_L1_run_cmp_tile_size_out_rsc_z;
  input [24:0] O_tiling_unit_L1_run_cmp_instr_bound_rsc_z;
  input [24:0] O_tiling_unit_L1_run_cmp_instr_tile_rsc_z;
  output O_tiling_unit_L1_run_cmp_ccs_ccore_start_rsc_dat;
  output O_tiling_unit_L1_run_cmp_ccs_ccore_en;


  // Interconnect Declarations
  wire run_wen;
  wire layer_instruction_in_rsci_wen_comp;
  wire [484:0] layer_instruction_in_rsci_idat_mxwt;
  wire O_instr_L1_out_rsci_wen_comp;
  wire O_instr_L2_out_rsci_wen_comp;
  wire O_instr_L3_out_rsci_wen_comp;
  wire I_instr_L1_out_rsci_wen_comp;
  wire I_instr_L2_out_rsci_wen_comp;
  wire I_instr_L3_out_rsci_wen_comp;
  wire W_instr_L1_out_rsci_wen_comp;
  wire W_instr_L2_out_rsci_wen_comp;
  wire W_instr_L3_out_rsci_wen_comp;
  reg ensig_cgo;
  reg ensig_cgo_1;
  reg ensig_cgo_2;
  reg ensig_cgo_3;
  reg ensig_cgo_4;
  reg [24:0] O_instr_L1_out_rsci_idat_49_25;
  reg [24:0] O_instr_L1_out_rsci_idat_24_0;
  reg [44:0] O_instr_L2_out_rsci_idat_89_45;
  reg [44:0] O_instr_L2_out_rsci_idat_44_0;
  reg [69:0] O_instr_L3_out_rsci_idat_139_70;
  reg [69:0] O_instr_L3_out_rsci_idat_69_0;
  reg [24:0] I_instr_L1_out_rsci_idat_49_25;
  reg [24:0] I_instr_L1_out_rsci_idat_24_0;
  reg [44:0] I_instr_L2_out_rsci_idat_89_45;
  reg [44:0] I_instr_L2_out_rsci_idat_44_0;
  reg [69:0] I_instr_L3_out_rsci_idat_139_70;
  reg [69:0] I_instr_L3_out_rsci_idat_69_0;
  reg [24:0] W_instr_L1_out_rsci_idat_49_25;
  reg [24:0] W_instr_L1_out_rsci_idat_24_0;
  reg [54:0] W_instr_L2_out_rsci_idat_109_55;
  reg [54:0] W_instr_L2_out_rsci_idat_54_0;
  reg [79:0] W_instr_L3_out_rsci_idat_159_80;
  reg [79:0] W_instr_L3_out_rsci_idat_79_0;
  wire [7:0] fsm_output;
  wire or_dcpl_1;
  wire or_dcpl_5;
  wire ensig_cgo_1_mx0;
  wire ensig_cgo_2_mx0;
  wire ensig_cgo_3_mx0;
  wire ensig_cgo_4_mx0;
  reg [484:0] layer_instruction_in_crt_sva;
  reg [4:0] O_tile_size_L1_sva;
  reg [4:0] I_tile_size_L1_sva;
  reg [4:0] W_tile_size_L1_sva;
  wire if_and_cse;
  wire if_and_2_cse;
  wire if_and_4_cse;
  wire if_and_10_cse;
  wire if_and_16_cse;
  reg reg_W_instr_L3_out_rsci_ivld_run_psct_cse;
  reg reg_W_instr_L2_out_rsci_ivld_run_psct_cse;
  reg reg_W_instr_L1_out_rsci_ivld_run_psct_cse;
  reg reg_I_instr_L1_out_rsci_ivld_run_psct_cse;
  reg reg_O_instr_L1_out_rsci_ivld_run_psct_cse;
  reg reg_layer_instruction_in_rsci_irdy_run_psct_cse;

  wire[4:0] if_mux_18_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [49:0] nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci_inst_O_instr_L1_out_rsci_idat;
  assign nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci_inst_O_instr_L1_out_rsci_idat
      = {O_instr_L1_out_rsci_idat_49_25 , O_instr_L1_out_rsci_idat_24_0};
  wire [89:0] nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci_inst_O_instr_L2_out_rsci_idat;
  assign nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci_inst_O_instr_L2_out_rsci_idat
      = {O_instr_L2_out_rsci_idat_89_45 , O_instr_L2_out_rsci_idat_44_0};
  wire [139:0] nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci_inst_O_instr_L3_out_rsci_idat;
  assign nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci_inst_O_instr_L3_out_rsci_idat
      = {O_instr_L3_out_rsci_idat_139_70 , O_instr_L3_out_rsci_idat_69_0};
  wire [49:0] nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci_inst_I_instr_L1_out_rsci_idat;
  assign nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci_inst_I_instr_L1_out_rsci_idat
      = {I_instr_L1_out_rsci_idat_49_25 , I_instr_L1_out_rsci_idat_24_0};
  wire [89:0] nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci_inst_I_instr_L2_out_rsci_idat;
  assign nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci_inst_I_instr_L2_out_rsci_idat
      = {I_instr_L2_out_rsci_idat_89_45 , I_instr_L2_out_rsci_idat_44_0};
  wire [139:0] nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci_inst_I_instr_L3_out_rsci_idat;
  assign nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci_inst_I_instr_L3_out_rsci_idat
      = {I_instr_L3_out_rsci_idat_139_70 , I_instr_L3_out_rsci_idat_69_0};
  wire [49:0] nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci_inst_W_instr_L1_out_rsci_idat;
  assign nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci_inst_W_instr_L1_out_rsci_idat
      = {W_instr_L1_out_rsci_idat_49_25 , W_instr_L1_out_rsci_idat_24_0};
  wire [109:0] nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci_inst_W_instr_L2_out_rsci_idat;
  assign nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci_inst_W_instr_L2_out_rsci_idat
      = {W_instr_L2_out_rsci_idat_109_55 , W_instr_L2_out_rsci_idat_54_0};
  wire [159:0] nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci_inst_W_instr_L3_out_rsci_idat;
  assign nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci_inst_W_instr_L3_out_rsci_idat
      = {W_instr_L3_out_rsci_idat_159_80 , W_instr_L3_out_rsci_idat_79_0};
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_layer_instruction_in_rsci
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_layer_instruction_in_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .layer_instruction_in_rsc_dat(layer_instruction_in_rsc_dat),
      .layer_instruction_in_rsc_vld(layer_instruction_in_rsc_vld),
      .layer_instruction_in_rsc_rdy(layer_instruction_in_rsc_rdy),
      .run_wen(run_wen),
      .layer_instruction_in_rsci_oswt(reg_layer_instruction_in_rsci_irdy_run_psct_cse),
      .layer_instruction_in_rsci_wen_comp(layer_instruction_in_rsci_wen_comp),
      .layer_instruction_in_rsci_idat_mxwt(layer_instruction_in_rsci_idat_mxwt)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .O_instr_L1_out_rsc_dat(O_instr_L1_out_rsc_dat),
      .O_instr_L1_out_rsc_vld(O_instr_L1_out_rsc_vld),
      .O_instr_L1_out_rsc_rdy(O_instr_L1_out_rsc_rdy),
      .run_wen(run_wen),
      .O_instr_L1_out_rsci_oswt(reg_O_instr_L1_out_rsci_ivld_run_psct_cse),
      .O_instr_L1_out_rsci_wen_comp(O_instr_L1_out_rsci_wen_comp),
      .O_instr_L1_out_rsci_idat(nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L1_out_rsci_inst_O_instr_L1_out_rsci_idat[49:0])
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .O_instr_L2_out_rsc_dat(O_instr_L2_out_rsc_dat),
      .O_instr_L2_out_rsc_vld(O_instr_L2_out_rsc_vld),
      .O_instr_L2_out_rsc_rdy(O_instr_L2_out_rsc_rdy),
      .run_wen(run_wen),
      .O_instr_L2_out_rsci_oswt(reg_W_instr_L1_out_rsci_ivld_run_psct_cse),
      .O_instr_L2_out_rsci_wen_comp(O_instr_L2_out_rsci_wen_comp),
      .O_instr_L2_out_rsci_idat(nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L2_out_rsci_inst_O_instr_L2_out_rsci_idat[89:0])
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .O_instr_L3_out_rsc_dat(O_instr_L3_out_rsc_dat),
      .O_instr_L3_out_rsc_vld(O_instr_L3_out_rsc_vld),
      .O_instr_L3_out_rsc_rdy(O_instr_L3_out_rsc_rdy),
      .run_wen(run_wen),
      .O_instr_L3_out_rsci_oswt(reg_W_instr_L2_out_rsci_ivld_run_psct_cse),
      .O_instr_L3_out_rsci_wen_comp(O_instr_L3_out_rsci_wen_comp),
      .O_instr_L3_out_rsci_idat(nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_O_instr_L3_out_rsci_inst_O_instr_L3_out_rsci_idat[139:0])
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .I_instr_L1_out_rsc_dat(I_instr_L1_out_rsc_dat),
      .I_instr_L1_out_rsc_vld(I_instr_L1_out_rsc_vld),
      .I_instr_L1_out_rsc_rdy(I_instr_L1_out_rsc_rdy),
      .run_wen(run_wen),
      .I_instr_L1_out_rsci_oswt(reg_I_instr_L1_out_rsci_ivld_run_psct_cse),
      .I_instr_L1_out_rsci_wen_comp(I_instr_L1_out_rsci_wen_comp),
      .I_instr_L1_out_rsci_idat(nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L1_out_rsci_inst_I_instr_L1_out_rsci_idat[49:0])
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .I_instr_L2_out_rsc_dat(I_instr_L2_out_rsc_dat),
      .I_instr_L2_out_rsc_vld(I_instr_L2_out_rsc_vld),
      .I_instr_L2_out_rsc_rdy(I_instr_L2_out_rsc_rdy),
      .run_wen(run_wen),
      .I_instr_L2_out_rsci_oswt(reg_W_instr_L2_out_rsci_ivld_run_psct_cse),
      .I_instr_L2_out_rsci_wen_comp(I_instr_L2_out_rsci_wen_comp),
      .I_instr_L2_out_rsci_idat(nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L2_out_rsci_inst_I_instr_L2_out_rsci_idat[89:0])
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .I_instr_L3_out_rsc_dat(I_instr_L3_out_rsc_dat),
      .I_instr_L3_out_rsc_vld(I_instr_L3_out_rsc_vld),
      .I_instr_L3_out_rsc_rdy(I_instr_L3_out_rsc_rdy),
      .run_wen(run_wen),
      .I_instr_L3_out_rsci_oswt(reg_W_instr_L3_out_rsci_ivld_run_psct_cse),
      .I_instr_L3_out_rsci_wen_comp(I_instr_L3_out_rsci_wen_comp),
      .I_instr_L3_out_rsci_idat(nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_I_instr_L3_out_rsci_inst_I_instr_L3_out_rsci_idat[139:0])
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .W_instr_L1_out_rsc_dat(W_instr_L1_out_rsc_dat),
      .W_instr_L1_out_rsc_vld(W_instr_L1_out_rsc_vld),
      .W_instr_L1_out_rsc_rdy(W_instr_L1_out_rsc_rdy),
      .run_wen(run_wen),
      .W_instr_L1_out_rsci_oswt(reg_W_instr_L1_out_rsci_ivld_run_psct_cse),
      .W_instr_L1_out_rsci_wen_comp(W_instr_L1_out_rsci_wen_comp),
      .W_instr_L1_out_rsci_idat(nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L1_out_rsci_inst_W_instr_L1_out_rsci_idat[49:0])
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .W_instr_L2_out_rsc_dat(W_instr_L2_out_rsc_dat),
      .W_instr_L2_out_rsc_vld(W_instr_L2_out_rsc_vld),
      .W_instr_L2_out_rsc_rdy(W_instr_L2_out_rsc_rdy),
      .run_wen(run_wen),
      .W_instr_L2_out_rsci_oswt(reg_W_instr_L2_out_rsci_ivld_run_psct_cse),
      .W_instr_L2_out_rsci_wen_comp(W_instr_L2_out_rsci_wen_comp),
      .W_instr_L2_out_rsci_idat(nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L2_out_rsci_inst_W_instr_L2_out_rsci_idat[109:0])
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .W_instr_L3_out_rsc_dat(W_instr_L3_out_rsc_dat),
      .W_instr_L3_out_rsc_vld(W_instr_L3_out_rsc_vld),
      .W_instr_L3_out_rsc_rdy(W_instr_L3_out_rsc_rdy),
      .run_wen(run_wen),
      .W_instr_L3_out_rsci_oswt(reg_W_instr_L3_out_rsci_ivld_run_psct_cse),
      .W_instr_L3_out_rsci_wen_comp(W_instr_L3_out_rsci_wen_comp),
      .W_instr_L3_out_rsci_idat(nl_config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_W_instr_L3_out_rsci_inst_W_instr_L3_out_rsci_idat[159:0])
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_wait_dp
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_wait_dp_inst
      (
      .ensig_cgo_iro(or_dcpl_5),
      .W_tiling_unit_L3_run_cmp_ccs_ccore_en(W_tiling_unit_L3_run_cmp_ccs_ccore_en),
      .ensig_cgo_iro_1(ensig_cgo_iro_1),
      .W_tiling_unit_L2_run_cmp_ccs_ccore_en(W_tiling_unit_L2_run_cmp_ccs_ccore_en),
      .ensig_cgo_iro_2(ensig_cgo_2_mx0),
      .O_tiling_unit_L3_run_cmp_ccs_ccore_en(O_tiling_unit_L3_run_cmp_ccs_ccore_en),
      .ensig_cgo_iro_3(ensig_cgo_3_mx0),
      .O_tiling_unit_L2_run_cmp_ccs_ccore_en(O_tiling_unit_L2_run_cmp_ccs_ccore_en),
      .ensig_cgo_iro_4(ensig_cgo_4_mx0),
      .O_tiling_unit_L1_run_cmp_ccs_ccore_en(O_tiling_unit_L1_run_cmp_ccs_ccore_en),
      .run_wen(run_wen),
      .ensig_cgo(ensig_cgo),
      .ensig_cgo_1(ensig_cgo_1),
      .ensig_cgo_2(ensig_cgo_2),
      .ensig_cgo_3(ensig_cgo_3),
      .ensig_cgo_4(ensig_cgo_4)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_staller
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_staller_inst
      (
      .run_wen(run_wen),
      .layer_instruction_in_rsci_wen_comp(layer_instruction_in_rsci_wen_comp),
      .O_instr_L1_out_rsci_wen_comp(O_instr_L1_out_rsci_wen_comp),
      .O_instr_L2_out_rsci_wen_comp(O_instr_L2_out_rsci_wen_comp),
      .O_instr_L3_out_rsci_wen_comp(O_instr_L3_out_rsci_wen_comp),
      .I_instr_L1_out_rsci_wen_comp(I_instr_L1_out_rsci_wen_comp),
      .I_instr_L2_out_rsci_wen_comp(I_instr_L2_out_rsci_wen_comp),
      .I_instr_L3_out_rsci_wen_comp(I_instr_L3_out_rsci_wen_comp),
      .W_instr_L1_out_rsci_wen_comp(W_instr_L1_out_rsci_wen_comp),
      .W_instr_L2_out_rsci_wen_comp(W_instr_L2_out_rsci_wen_comp),
      .W_instr_L3_out_rsci_wen_comp(W_instr_L3_out_rsci_wen_comp)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_run_fsm
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_run_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign if_and_cse = run_wen & (fsm_output[6]);
  assign if_and_2_cse = run_wen & (fsm_output[5]);
  assign if_and_4_cse = run_wen & (fsm_output[4]);
  assign if_and_10_cse = run_wen & (fsm_output[3]);
  assign if_and_16_cse = run_wen & (fsm_output[2]);
  assign ensig_cgo_4_mx0 = or_dcpl_1 | (fsm_output[1]) | (fsm_output[4]);
  assign ensig_cgo_3_mx0 = (fsm_output[5:3]!=3'b000);
  assign ensig_cgo_2_mx0 = or_dcpl_5 | (fsm_output[4]);
  assign ensig_cgo_1_mx0 = (fsm_output[5:4]!=2'b00);
  assign or_dcpl_1 = (fsm_output[3:2]!=2'b00);
  assign or_dcpl_5 = (fsm_output[6:5]!=2'b00);
  assign W_tiling_unit_L3_run_cmp_loops_bound_rsc_dat = layer_instruction_in_crt_sva[389:310];
  assign W_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat = layer_instruction_in_crt_sva[394:390];
  assign W_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat = {5'b0, W_tiling_unit_L2_run_cmp_tile_size_out_rsc_z};
  assign W_tiling_unit_L3_run_cmp_ccs_ccore_start_rsc_dat = fsm_output[5];
  assign W_tiling_unit_L2_run_cmp_loops_bound_rsc_dat = layer_instruction_in_crt_sva[449:395];
  assign W_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat = layer_instruction_in_crt_sva[454:450];
  assign W_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat = {6'b0, O_tiling_unit_L1_run_cmp_tile_size_out_rsc_z};
  assign W_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat = fsm_output[4];
  assign O_tiling_unit_L3_run_cmp_loops_bound_rsc_dat = MUX_v_70_2_2((layer_instruction_in_crt_sva[69:0]),
      (layer_instruction_in_crt_sva[224:155]), fsm_output[5]);
  assign O_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat = MUX_v_5_2_2((layer_instruction_in_crt_sva[74:70]),
      (layer_instruction_in_crt_sva[229:225]), fsm_output[5]);
  assign O_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat = {5'b0, O_tiling_unit_L2_run_cmp_tile_size_out_rsc_z};
  assign O_tiling_unit_L2_run_cmp_loops_bound_rsc_dat = MUX_v_45_2_2((layer_instruction_in_crt_sva[119:75]),
      (layer_instruction_in_crt_sva[274:230]), fsm_output[4]);
  assign O_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat = MUX_v_5_2_2((layer_instruction_in_crt_sva[124:120]),
      (layer_instruction_in_crt_sva[279:275]), fsm_output[4]);
  assign if_mux_18_nl = MUX_v_5_2_2(O_tile_size_L1_sva, I_tile_size_L1_sva, fsm_output[4]);
  assign O_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat = {4'b0, if_mux_18_nl};
  assign O_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat = (fsm_output[4:3]!=2'b00);
  assign O_tiling_unit_L1_run_cmp_loops_bound_rsc_dat = MUX1HOT_v_25_3_2((layer_instruction_in_rsci_idat_mxwt[149:125]),
      (layer_instruction_in_crt_sva[304:280]), (layer_instruction_in_crt_sva[479:455]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
  assign O_tiling_unit_L1_run_cmp_loops_relevancy_rsc_dat = MUX1HOT_v_5_3_2((layer_instruction_in_rsci_idat_mxwt[154:150]),
      (layer_instruction_in_crt_sva[309:305]), (layer_instruction_in_crt_sva[484:480]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
  assign O_tiling_unit_L1_run_cmp_tile_size_in_rsc_dat = MUX1HOT_v_5_3_2(O_tile_size_L1_sva,
      I_tile_size_L1_sva, W_tile_size_L1_sva, {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3])});
  assign O_tiling_unit_L1_run_cmp_ccs_ccore_start_rsc_dat = or_dcpl_1 | (fsm_output[1]);
  assign CGHpart_irsig_1 = ensig_cgo_1_mx0;
  always @(posedge clk) begin
    if ( rst ) begin
      W_instr_L3_out_rsci_idat_79_0 <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
      W_instr_L3_out_rsci_idat_159_80 <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
      I_instr_L3_out_rsci_idat_69_0 <= 70'b0000000000000000000000000000000000000000000000000000000000000000000000;
      I_instr_L3_out_rsci_idat_139_70 <= 70'b0000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( if_and_cse ) begin
      W_instr_L3_out_rsci_idat_79_0 <= W_tiling_unit_L3_run_cmp_instr_bound_rsc_z;
      W_instr_L3_out_rsci_idat_159_80 <= W_tiling_unit_L3_run_cmp_instr_tile_rsc_z;
      I_instr_L3_out_rsci_idat_69_0 <= O_tiling_unit_L3_run_cmp_instr_bound_rsc_z;
      I_instr_L3_out_rsci_idat_139_70 <= O_tiling_unit_L3_run_cmp_instr_tile_rsc_z;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_instr_L2_out_rsci_idat_54_0 <= 55'b0000000000000000000000000000000000000000000000000000000;
      W_instr_L2_out_rsci_idat_109_55 <= 55'b0000000000000000000000000000000000000000000000000000000;
      I_instr_L2_out_rsci_idat_44_0 <= 45'b000000000000000000000000000000000000000000000;
      I_instr_L2_out_rsci_idat_89_45 <= 45'b000000000000000000000000000000000000000000000;
      O_instr_L3_out_rsci_idat_69_0 <= 70'b0000000000000000000000000000000000000000000000000000000000000000000000;
      O_instr_L3_out_rsci_idat_139_70 <= 70'b0000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( if_and_2_cse ) begin
      W_instr_L2_out_rsci_idat_54_0 <= W_tiling_unit_L2_run_cmp_instr_bound_rsc_z;
      W_instr_L2_out_rsci_idat_109_55 <= W_tiling_unit_L2_run_cmp_instr_tile_rsc_z;
      I_instr_L2_out_rsci_idat_44_0 <= O_tiling_unit_L2_run_cmp_instr_bound_rsc_z;
      I_instr_L2_out_rsci_idat_89_45 <= O_tiling_unit_L2_run_cmp_instr_tile_rsc_z;
      O_instr_L3_out_rsci_idat_69_0 <= O_tiling_unit_L3_run_cmp_instr_bound_rsc_z;
      O_instr_L3_out_rsci_idat_139_70 <= O_tiling_unit_L3_run_cmp_instr_tile_rsc_z;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_instr_L1_out_rsci_idat_24_0 <= 25'b0000000000000000000000000;
      W_instr_L1_out_rsci_idat_49_25 <= 25'b0000000000000000000000000;
      O_instr_L2_out_rsci_idat_44_0 <= 45'b000000000000000000000000000000000000000000000;
      O_instr_L2_out_rsci_idat_89_45 <= 45'b000000000000000000000000000000000000000000000;
      W_tile_size_L1_sva <= 5'b00001;
    end
    else if ( if_and_4_cse ) begin
      W_instr_L1_out_rsci_idat_24_0 <= O_tiling_unit_L1_run_cmp_instr_bound_rsc_z;
      W_instr_L1_out_rsci_idat_49_25 <= O_tiling_unit_L1_run_cmp_instr_tile_rsc_z;
      O_instr_L2_out_rsci_idat_44_0 <= O_tiling_unit_L2_run_cmp_instr_bound_rsc_z;
      O_instr_L2_out_rsci_idat_89_45 <= O_tiling_unit_L2_run_cmp_instr_tile_rsc_z;
      W_tile_size_L1_sva <= O_tiling_unit_L1_run_cmp_tile_size_out_rsc_z;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_instr_L1_out_rsci_idat_24_0 <= 25'b0000000000000000000000000;
      I_instr_L1_out_rsci_idat_49_25 <= 25'b0000000000000000000000000;
      I_tile_size_L1_sva <= 5'b00001;
    end
    else if ( if_and_10_cse ) begin
      I_instr_L1_out_rsci_idat_24_0 <= O_tiling_unit_L1_run_cmp_instr_bound_rsc_z;
      I_instr_L1_out_rsci_idat_49_25 <= O_tiling_unit_L1_run_cmp_instr_tile_rsc_z;
      I_tile_size_L1_sva <= O_tiling_unit_L1_run_cmp_tile_size_out_rsc_z;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_instr_L1_out_rsci_idat_24_0 <= 25'b0000000000000000000000000;
      O_instr_L1_out_rsci_idat_49_25 <= 25'b0000000000000000000000000;
      O_tile_size_L1_sva <= 5'b00001;
    end
    else if ( if_and_16_cse ) begin
      O_instr_L1_out_rsci_idat_24_0 <= O_tiling_unit_L1_run_cmp_instr_bound_rsc_z;
      O_instr_L1_out_rsci_idat_49_25 <= O_tiling_unit_L1_run_cmp_instr_tile_rsc_z;
      O_tile_size_L1_sva <= O_tiling_unit_L1_run_cmp_tile_size_out_rsc_z;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ensig_cgo_4 <= 1'b0;
      ensig_cgo_3 <= 1'b0;
      ensig_cgo_2 <= 1'b0;
      ensig_cgo_1 <= 1'b0;
      ensig_cgo <= 1'b0;
      reg_W_instr_L3_out_rsci_ivld_run_psct_cse <= 1'b0;
      reg_W_instr_L2_out_rsci_ivld_run_psct_cse <= 1'b0;
      reg_W_instr_L1_out_rsci_ivld_run_psct_cse <= 1'b0;
      reg_I_instr_L1_out_rsci_ivld_run_psct_cse <= 1'b0;
      reg_O_instr_L1_out_rsci_ivld_run_psct_cse <= 1'b0;
      reg_layer_instruction_in_rsci_irdy_run_psct_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      ensig_cgo_4 <= ensig_cgo_4_mx0;
      ensig_cgo_3 <= ensig_cgo_3_mx0;
      ensig_cgo_2 <= ensig_cgo_2_mx0;
      ensig_cgo_1 <= ensig_cgo_1_mx0;
      ensig_cgo <= or_dcpl_5;
      reg_W_instr_L3_out_rsci_ivld_run_psct_cse <= fsm_output[6];
      reg_W_instr_L2_out_rsci_ivld_run_psct_cse <= fsm_output[5];
      reg_W_instr_L1_out_rsci_ivld_run_psct_cse <= fsm_output[4];
      reg_I_instr_L1_out_rsci_ivld_run_psct_cse <= fsm_output[3];
      reg_O_instr_L1_out_rsci_ivld_run_psct_cse <= fsm_output[2];
      reg_layer_instruction_in_rsci_irdy_run_psct_cse <= (fsm_output[7]) | (fsm_output[0]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer_instruction_in_crt_sva <= 485'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      layer_instruction_in_crt_sva <= layer_instruction_in_rsci_idat_mxwt;
    end
  end

  function automatic [24:0] MUX1HOT_v_25_3_2;
    input [24:0] input_2;
    input [24:0] input_1;
    input [24:0] input_0;
    input [2:0] sel;
    reg [24:0] result;
  begin
    result = input_0 & {25{sel[0]}};
    result = result | ( input_1 & {25{sel[1]}});
    result = result | ( input_2 & {25{sel[2]}});
    MUX1HOT_v_25_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [44:0] MUX_v_45_2_2;
    input [44:0] input_0;
    input [44:0] input_1;
    input [0:0] sel;
    reg [44:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_45_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [69:0] MUX_v_70_2_2;
    input [69:0] input_0;
    input [69:0] input_1;
    input [0:0] sel;
    reg [69:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_70_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run
    (
  clk, rst, O_wr_data_rsc_dat, O_wr_data_rsc_vld, O_wr_data_rsc_rdy, O_rd_data_rsc_dat,
      O_rd_data_rsc_vld, O_rd_data_rsc_rdy, I_wr_data_rsc_dat, I_wr_data_rsc_vld,
      I_wr_data_rsc_rdy, W_wr_data_rsc_dat, W_wr_data_rsc_vld, W_wr_data_rsc_rdy,
      wr_data_zero_guard_rsc_dat, wr_data_zero_guard_rsc_vld, wr_data_zero_guard_rsc_rdy,
      O_instr_in_rsc_dat, O_instr_in_rsc_vld, O_instr_in_rsc_rdy, I_instr_in_rsc_dat,
      I_instr_in_rsc_vld, I_instr_in_rsc_rdy, W_instr_in_rsc_dat, W_instr_in_rsc_vld,
      W_instr_in_rsc_rdy
);
  input clk;
  input rst;
  input [15:0] O_wr_data_rsc_dat;
  input O_wr_data_rsc_vld;
  output O_wr_data_rsc_rdy;
  output [15:0] O_rd_data_rsc_dat;
  output O_rd_data_rsc_vld;
  input O_rd_data_rsc_rdy;
  input [15:0] I_wr_data_rsc_dat;
  input I_wr_data_rsc_vld;
  output I_wr_data_rsc_rdy;
  input [15:0] W_wr_data_rsc_dat;
  input W_wr_data_rsc_vld;
  output W_wr_data_rsc_rdy;
  input wr_data_zero_guard_rsc_dat;
  input wr_data_zero_guard_rsc_vld;
  output wr_data_zero_guard_rsc_rdy;
  input [49:0] O_instr_in_rsc_dat;
  input O_instr_in_rsc_vld;
  output O_instr_in_rsc_rdy;
  input [49:0] I_instr_in_rsc_dat;
  input I_instr_in_rsc_vld;
  output I_instr_in_rsc_rdy;
  input [49:0] W_instr_in_rsc_dat;
  input W_instr_in_rsc_vld;
  output W_instr_in_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire O_wr_data_rsci_ivld_mxwt;
  wire [15:0] O_wr_data_rsci_idat_mxwt;
  wire O_rd_data_rsci_irdy_mxwt;
  reg [15:0] O_rd_data_rsci_idat;
  wire I_wr_data_rsci_ivld_mxwt;
  wire [15:0] I_wr_data_rsci_idat_mxwt;
  wire W_wr_data_rsci_ivld_mxwt;
  wire [15:0] W_wr_data_rsci_idat_mxwt;
  wire wr_data_zero_guard_rsci_ivld_mxwt;
  wire wr_data_zero_guard_rsci_idat_mxwt;
  wire O_instr_in_rsci_wen_comp;
  wire [49:0] O_instr_in_rsci_idat_mxwt;
  wire I_instr_in_rsci_wen_comp;
  wire [49:0] I_instr_in_rsci_idat_mxwt;
  wire W_instr_in_rsci_wen_comp;
  wire [49:0] W_instr_in_rsci_idat_mxwt;
  wire [1:0] fsm_output;
  wire [1:0] mux1h_1_tmp;
  wire aif_7_equal_tmp;
  wire [1:0] mux_188_tmp;
  wire if_6_aif_equal_tmp;
  wire [4:0] if_6_if_3_acc_tmp;
  wire [5:0] nl_if_6_if_3_acc_tmp;
  wire [4:0] if_6_if_1_acc_tmp;
  wire [5:0] nl_if_6_if_1_acc_tmp;
  wire [4:0] if_6_if_6_mux1h_tmp;
  wire if_6_else_if_equal_tmp;
  wire aif_equal_tmp;
  wire oif_2_unequal_tmp;
  wire oif_1_unequal_tmp;
  wire oif_unequal_tmp;
  wire if_for_if_for_and_26_tmp;
  wire if_for_if_for_and_28_tmp;
  wire if_for_if_for_and_27_tmp;
  wire if_5_else_or_tmp_2;
  wire if_10_if_equal_1_tmp;
  wire if_9_if_equal_1_tmp;
  wire [1:0] mux1h_7_tmp;
  wire or_tmp_2;
  wire and_tmp;
  wire and_tmp_1;
  wire or_tmp_5;
  wire mux_tmp_4;
  wire mux_tmp_6;
  wire or_tmp_10;
  wire mux_tmp_11;
  wire and_dcpl;
  wire and_tmp_14;
  wire mux_tmp_14;
  wire nor_tmp_8;
  wire not_tmp_8;
  wire not_tmp_9;
  wire mux_tmp_24;
  wire not_tmp_14;
  wire not_tmp_15;
  wire mux_tmp_34;
  wire or_tmp_51;
  wire nor_tmp_25;
  wire and_tmp_40;
  wire nor_tmp_26;
  wire or_dcpl_11;
  wire not_tmp_25;
  wire or_tmp_73;
  wire or_dcpl_14;
  wire nor_tmp_39;
  wire nor_tmp_43;
  wire or_tmp_93;
  wire mux_tmp_67;
  wire or_tmp_96;
  wire or_tmp_97;
  wire or_tmp_98;
  wire and_dcpl_19;
  wire or_dcpl_19;
  wire or_dcpl_21;
  wire or_dcpl_22;
  wire or_dcpl_23;
  wire or_dcpl_25;
  wire or_dcpl_27;
  wire or_dcpl_28;
  wire or_dcpl_29;
  wire or_dcpl_31;
  wire or_dcpl_32;
  wire or_dcpl_33;
  wire or_dcpl_34;
  wire or_dcpl_35;
  wire or_dcpl_36;
  wire or_dcpl_37;
  wire or_dcpl_38;
  wire or_dcpl_39;
  wire or_dcpl_40;
  wire or_dcpl_41;
  wire or_dcpl_43;
  wire or_dcpl_44;
  wire or_dcpl_45;
  wire or_dcpl_47;
  wire or_dcpl_48;
  wire or_dcpl_49;
  wire or_dcpl_50;
  wire or_dcpl_51;
  wire or_dcpl_52;
  wire or_dcpl_53;
  wire or_dcpl_54;
  wire or_dcpl_55;
  wire or_dcpl_56;
  wire or_dcpl_57;
  wire or_dcpl_58;
  wire or_dcpl_59;
  wire or_dcpl_60;
  wire or_dcpl_61;
  wire or_dcpl_62;
  wire or_dcpl_63;
  wire or_dcpl_64;
  wire or_dcpl_65;
  wire or_dcpl_66;
  wire or_dcpl_67;
  wire or_dcpl_68;
  wire or_dcpl_69;
  wire or_dcpl_70;
  wire or_dcpl_71;
  wire or_dcpl_72;
  wire or_dcpl_73;
  wire not_tmp_47;
  wire mux_tmp_76;
  wire or_dcpl_78;
  wire or_dcpl_80;
  wire or_dcpl_81;
  wire or_dcpl_82;
  wire or_dcpl_84;
  wire or_dcpl_87;
  wire or_dcpl_88;
  wire or_dcpl_89;
  wire or_dcpl_90;
  wire or_dcpl_91;
  wire or_dcpl_92;
  wire or_dcpl_94;
  wire or_dcpl_95;
  wire or_dcpl_97;
  wire or_dcpl_98;
  wire or_dcpl_99;
  wire or_dcpl_100;
  wire or_dcpl_101;
  wire or_dcpl_102;
  wire or_dcpl_103;
  wire or_dcpl_104;
  wire or_dcpl_105;
  wire or_dcpl_106;
  wire or_dcpl_107;
  wire or_dcpl_108;
  wire or_dcpl_109;
  wire or_dcpl_110;
  wire or_dcpl_111;
  wire or_dcpl_112;
  wire or_dcpl_113;
  wire or_dcpl_114;
  wire or_dcpl_115;
  wire or_dcpl_116;
  wire or_dcpl_117;
  wire or_dcpl_118;
  wire or_dcpl_119;
  wire or_dcpl_120;
  wire or_dcpl_121;
  wire or_dcpl_122;
  wire or_dcpl_123;
  wire or_dcpl_124;
  wire or_dcpl_125;
  wire or_dcpl_126;
  wire or_dcpl_127;
  wire or_dcpl_128;
  wire or_dcpl_129;
  wire or_dcpl_130;
  wire or_dcpl_131;
  wire or_dcpl_132;
  wire and_tmp_56;
  wire or_tmp_105;
  wire mux_tmp_77;
  wire or_tmp_106;
  wire mux_tmp_78;
  wire and_tmp_57;
  wire mux_tmp_79;
  wire not_tmp_56;
  wire mux_tmp_84;
  wire or_dcpl_136;
  wire or_dcpl_137;
  wire or_dcpl_138;
  wire or_dcpl_139;
  wire nor_tmp_65;
  wire mux_tmp_89;
  wire mux_tmp_91;
  wire or_dcpl_142;
  wire or_dcpl_143;
  wire or_dcpl_146;
  wire or_dcpl_147;
  wire or_dcpl_150;
  wire or_dcpl_151;
  wire or_dcpl_154;
  wire or_dcpl_155;
  wire or_dcpl_158;
  wire or_dcpl_161;
  wire or_dcpl_164;
  wire or_dcpl_167;
  wire or_dcpl_168;
  wire or_dcpl_171;
  wire or_dcpl_174;
  wire or_dcpl_177;
  wire or_dcpl_180;
  wire or_dcpl_181;
  wire or_dcpl_184;
  wire or_dcpl_187;
  wire or_dcpl_190;
  wire or_dcpl_193;
  wire or_dcpl_226;
  wire mux_tmp_94;
  wire mux_tmp_96;
  wire mux_tmp_98;
  wire or_dcpl_237;
  wire or_tmp_143;
  wire mux_tmp_113;
  wire or_tmp_162;
  wire not_tmp_93;
  wire mux_tmp_129;
  wire nand_tmp_25;
  wire nand_tmp_27;
  wire mux_tmp_134;
  wire or_tmp_171;
  wire nand_tmp_28;
  wire nor_tmp_110;
  wire mux_tmp_143;
  wire nand_tmp_29;
  wire mux_tmp_144;
  wire nand_tmp_30;
  wire mux_tmp_153;
  wire nand_tmp_31;
  wire nand_tmp_32;
  wire mux_tmp_161;
  wire nand_tmp_33;
  wire mux_tmp_170;
  wire nand_tmp_34;
  wire mux_tmp_171;
  wire nand_tmp_35;
  wire mux_tmp_180;
  wire or_tmp_200;
  wire mux_tmp_189;
  wire and_tmp_80;
  wire or_tmp_204;
  wire mux_tmp_202;
  wire and_tmp_81;
  wire or_dcpl_246;
  wire or_dcpl_248;
  wire and_tmp_93;
  wire mux_tmp_224;
  wire mux_tmp_226;
  wire mux_tmp_231;
  wire mux_tmp_232;
  wire and_tmp_98;
  wire and_dcpl_28;
  wire or_tmp_242;
  wire land_8_lpi_1_dfm_1;
  wire skid_buf_wr_zero_guard_peek_slc_skid_buf_wr_zero_guard_regs_skid_buf_wr_zero_guard_rd_ptr_1_0_cse_sva_mx0;
  wire O_data_vld_sva_dfm_4_mx0;
  wire W_data_vld_sva_mx0;
  wire if_6_unequal_tmp_2;
  wire I_data_vld_sva_mx0;
  wire if_6_unequal_tmp_3;
  reg O_data_vld_sva;
  wire O_write_flag_sva_mx0;
  wire land_lpi_1_dfm_1;
  wire [4:0] W_irrel_cnt_sva_dfm_mx0;
  wire [4:0] I_irrel_cnt_sva_dfm_mx0;
  wire skid_buf_top_rd_ptr_sva_1_mx1;
  wire skid_buf_top_rd_ptr_sva_0_mx1;
  wire skid_buf_top_wr_ptr_sva_0_mx1;
  wire skid_buf_top_wr_ptr_sva_1_mx1;
  wire land_5_lpi_1_dfm_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1;
  wire land_2_lpi_1_dfm_2;
  wire lor_4_lpi_1_dfm_1;
  wire O_mac_irrel_at_max_sva_dfm_mx0;
  reg flags_top_1_1_sva;
  wire lor_2_lpi_1_dfm_1;
  wire aif_3_land_lpi_1_dfm_mx0;
  wire lor_3_lpi_1_dfm_1;
  wire lor_1_lpi_1_dfm_1;
  wire aif_2_land_1_lpi_1_dfm_mx0;
  reg data_zg_sva;
  wire W_write_flag_sva_mx0;
  reg W_data_vld_sva_dfm_1_1;
  wire I_write_flag_sva_mx0;
  reg I_data_vld_sva_dfm_1_1;
  reg skid_buf_top_rd_ptr_sva_1;
  reg skid_buf_top_rd_ptr_sva_0;
  wire if_5_if_nbw_stat_sva_mx1;
  wire and_17_m1c_1;
  wire and_16_m1c_1;
  reg or_svs_1;
  reg skid_buf_top_wr_ptr_sva_1;
  wire skid_buf_top_push_1_xor_psp_1;
  wire skid_buf_top_push_1_skid_buf_top_push_1_nand_seb_1;
  reg skid_buf_top_wr_ptr_sva_dfm_1_1;
  reg skid_buf_top_wr_ptr_sva_0;
  reg skid_buf_top_push_nor_psp;
  reg [49:0] W_instr_in_crt_lpi_1_dfm_1;
  reg [49:0] I_instr_in_crt_lpi_1_dfm_1;
  reg operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1_1;
  reg if_5_and_svs_1;
  wire skid_buf_top_pop_1_xor_psp_1;
  wire else_8_land_lpi_1_dfm_mx1;
  wire land_9_lpi_1_dfm_1;
  reg skid_buf_wr_zero_guard_wr_ptr_sva;
  reg [1:0] skid_buf_top_cnt_sva;
  reg main_stage_0_2;
  reg mux_124_itm_1;
  reg land_9_lpi_1_dfm_1_1;
  reg O_mac_irrel_at_max_sva;
  reg [3:0] W_irrel_cnt_sva_4_1;
  reg W_irrel_cnt_sva_0;
  reg W_mac_irrel_at_maxBuf_sva;
  reg [3:0] I_irrel_cnt_sva_4_1;
  reg I_irrel_cnt_sva_0;
  reg I_mac_irrel_at_maxBuf_sva;
  reg skid_buf_wr_zero_guard_rd_ptr_sva;
  reg [4:0] W_wr_pntr_sva;
  reg [4:0] I_wr_pntr_sva;
  reg [4:0] O_mac_pntr_sva;
  reg skid_buf_top_push_and_psp;
  reg skid_buf_top_push_and_1_psp;
  reg skid_buf_wr_zero_guard_regs_0_sva_dfm_1;
  reg skid_buf_wr_zero_guard_regs_1_sva_dfm_1;
  reg flags_wr_zero_guard_sva;
  wire [4:0] if_10_if_ac_int_cctor_sva_1;
  wire [5:0] nl_if_10_if_ac_int_cctor_sva_1;
  wire [4:0] if_9_if_ac_int_cctor_sva_1;
  wire [5:0] nl_if_9_if_ac_int_cctor_sva_1;
  wire [1:0] skid_buf_top_cnt_sva_mx1;
  wire skid_buf_top_pop_1_skid_buf_top_pop_1_nand_seb_1;
  wire nand_11_ssc_1;
  wire and_47_ssc_1;
  wire or_360_tmp;
  wire skid_buf_top_peek_and_m1c;
  wire or_364_tmp;
  wire skid_buf_top_peek_and_4_m1c;
  wire or_368_tmp;
  wire skid_buf_top_peek_and_5_m1c;
  wire if_5_if_and_3_m1c;
  wire if_5_if_and_4_m1c;
  wire if_5_if_and_5_m1c;
  reg reg_wr_data_zero_guard_rsci_oswt_cse;
  reg reg_W_wr_data_rsci_irdy_run_psct_cse;
  reg reg_I_wr_data_rsci_irdy_run_psct_cse;
  reg reg_O_rd_data_rsci_ivld_run_psct_cse;
  reg reg_O_wr_data_rsci_irdy_run_psct_cse;
  wire W_mac_pntr_and_cse;
  wire flags_wr_zero_guard_and_cse;
  wire nor_108_cse;
  wire W_mac_irrel_at_maxBuf_and_cse;
  wire skid_buf_top_push_and_2_cse;
  wire operator_2_false_5_operator_2_false_5_operator_2_false_5_or_cse;
  wire or_570_cse;
  wire mux_420_cse;
  wire [1:0] mux_124_cse;
  wire or_1_cse;
  wire or_558_cse;
  wire and_295_cse;
  wire or_18_cse;
  wire or_569_cse;
  wire nor_110_cse;
  wire or_359_cse;
  wire or_363_cse;
  wire or_367_cse;
  wire mux_554_cse;
  wire and_306_cse;
  wire mux_396_cse;
  wire or_557_cse;
  wire mux_342_cse;
  wire nand_78_cse;
  wire mux_343_cse;
  wire mux_346_cse;
  wire or_399_cse;
  wire or_400_cse;
  wire or_401_cse;
  wire mux_405_cse;
  wire mux_460_cse;
  wire else_3_land_lpi_1_dfm_mx0w0;
  reg else_3_land_lpi_1_dfm;
  wire [4:0] if_6_if_if_6_if_and_1_itm;
  wire if_6_or_itm;
  wire mux_426_itm;
  wire mux_571_itm;
  wire [15:0] z_out_2;
  wire [31:0] nl_z_out_2;
  wire [1:0] z_out_3;
  wire [2:0] nl_z_out_3;
  reg [4:0] O_mac_tile_bound_0_lpi_1;
  reg [4:0] I_mac_tile_bound_0_lpi_1;
  reg [4:0] W_mac_tile_bound_0_lpi_1;
  reg [4:0] O_mac_tile_bound_1_lpi_1;
  reg [4:0] I_mac_tile_bound_1_lpi_1;
  reg [4:0] W_mac_tile_bound_1_lpi_1;
  reg [4:0] O_mac_tile_bound_2_lpi_1;
  reg [4:0] I_mac_tile_bound_2_lpi_1;
  reg [4:0] W_mac_tile_bound_2_lpi_1;
  reg [4:0] O_mac_tile_bound_3_lpi_1;
  reg [4:0] I_mac_tile_bound_3_lpi_1;
  reg [4:0] W_mac_tile_bound_3_lpi_1;
  reg [4:0] O_mac_tile_bound_4_lpi_1;
  reg [4:0] I_mac_tile_bound_4_lpi_1;
  reg [4:0] W_mac_tile_bound_4_lpi_1;
  reg [15:0] skid_buf_top_regs_data_1_0_sva;
  reg [15:0] skid_buf_top_regs_data_0_0_sva;
  reg [15:0] skid_buf_top_regs_data_2_0_sva;
  reg [1:0] skid_buf_wr_zero_guard_cnt_sva;
  reg [15:0] O_mem_15_sva;
  reg [15:0] O_mem_16_sva;
  reg [15:0] O_mem_14_sva;
  reg [15:0] O_mem_17_sva;
  reg [15:0] O_mem_13_sva;
  reg [15:0] O_mem_18_sva;
  reg [15:0] O_mem_12_sva;
  reg [15:0] O_mem_19_sva;
  reg [15:0] O_mem_11_sva;
  reg [15:0] O_mem_20_sva;
  reg [15:0] O_mem_10_sva;
  reg [15:0] O_mem_21_sva;
  reg [15:0] O_mem_9_sva;
  reg [15:0] O_mem_22_sva;
  reg [15:0] O_mem_8_sva;
  reg [15:0] O_mem_23_sva;
  reg [15:0] O_mem_7_sva;
  reg [15:0] O_mem_24_sva;
  reg [15:0] O_mem_6_sva;
  reg [15:0] O_mem_25_sva;
  reg [15:0] O_mem_5_sva;
  reg [15:0] O_mem_26_sva;
  reg [15:0] O_mem_4_sva;
  reg [15:0] O_mem_27_sva;
  reg [15:0] O_mem_3_sva;
  reg [15:0] O_mem_28_sva;
  reg [15:0] O_mem_2_sva;
  reg [15:0] O_mem_29_sva;
  reg [15:0] O_mem_1_sva;
  reg [15:0] O_mem_30_sva;
  reg [15:0] O_mem_0_sva;
  reg [15:0] O_mem_31_sva;
  reg [15:0] O_write_data_data_sva;
  reg [4:0] O_vld_zg_pntr_sva;
  reg [15:0] I_mem_15_sva;
  reg [15:0] I_mem_16_sva;
  reg [15:0] I_mem_14_sva;
  reg [15:0] I_mem_17_sva;
  reg [15:0] I_mem_13_sva;
  reg [15:0] I_mem_18_sva;
  reg [15:0] I_mem_12_sva;
  reg [15:0] I_mem_19_sva;
  reg [15:0] I_mem_11_sva;
  reg [15:0] I_mem_20_sva;
  reg [15:0] I_mem_10_sva;
  reg [15:0] I_mem_21_sva;
  reg [15:0] I_mem_9_sva;
  reg [15:0] I_mem_22_sva;
  reg [15:0] I_mem_8_sva;
  reg [15:0] I_mem_23_sva;
  reg [15:0] I_mem_7_sva;
  reg [15:0] I_mem_24_sva;
  reg [15:0] I_mem_6_sva;
  reg [15:0] I_mem_25_sva;
  reg [15:0] I_mem_5_sva;
  reg [15:0] I_mem_26_sva;
  reg [15:0] I_mem_4_sva;
  reg [15:0] I_mem_27_sva;
  reg [15:0] I_mem_3_sva;
  reg [15:0] I_mem_28_sva;
  reg [15:0] I_mem_2_sva;
  reg [15:0] I_mem_29_sva;
  reg [15:0] I_mem_1_sva;
  reg [15:0] I_mem_30_sva;
  reg [15:0] I_mem_0_sva;
  reg [15:0] I_mem_31_sva;
  reg [4:0] I_mac_pntr_sva;
  reg [15:0] W_mem_15_sva;
  reg [15:0] W_mem_16_sva;
  reg [15:0] W_mem_14_sva;
  reg [15:0] W_mem_17_sva;
  reg [15:0] W_mem_13_sva;
  reg [15:0] W_mem_18_sva;
  reg [15:0] W_mem_12_sva;
  reg [15:0] W_mem_19_sva;
  reg [15:0] W_mem_11_sva;
  reg [15:0] W_mem_20_sva;
  reg [15:0] W_mem_10_sva;
  reg [15:0] W_mem_21_sva;
  reg [15:0] W_mem_9_sva;
  reg [15:0] W_mem_22_sva;
  reg [15:0] W_mem_8_sva;
  reg [15:0] W_mem_23_sva;
  reg [15:0] W_mem_7_sva;
  reg [15:0] W_mem_24_sva;
  reg [15:0] W_mem_6_sva;
  reg [15:0] W_mem_25_sva;
  reg [15:0] W_mem_5_sva;
  reg [15:0] W_mem_26_sva;
  reg [15:0] W_mem_4_sva;
  reg [15:0] W_mem_27_sva;
  reg [15:0] W_mem_3_sva;
  reg [15:0] W_mem_28_sva;
  reg [15:0] W_mem_2_sva;
  reg [15:0] W_mem_29_sva;
  reg [15:0] W_mem_1_sva;
  reg [15:0] W_mem_30_sva;
  reg [15:0] W_mem_0_sva;
  reg [15:0] W_mem_31_sva;
  reg [4:0] W_mac_pntr_sva;
  reg [4:0] O_mac_counter_2_sva;
  reg [4:0] O_mac_counter_1_sva;
  reg [4:0] O_mac_counter_3_sva;
  reg [4:0] O_mac_counter_0_sva;
  reg [4:0] O_mac_counter_4_sva;
  reg [4:0] I_mac_counter_2_sva;
  reg [4:0] I_mac_counter_1_sva;
  reg [4:0] I_mac_counter_3_sva;
  reg [4:0] I_mac_counter_0_sva;
  reg [4:0] I_mac_counter_4_sva;
  reg [4:0] W_mac_counter_2_sva;
  reg [4:0] W_mac_counter_1_sva;
  reg [4:0] W_mac_counter_3_sva;
  reg [4:0] W_mac_counter_0_sva;
  reg [4:0] W_mac_counter_4_sva;
  reg [49:0] O_instr_in_crt_lpi_1_dfm;
  reg aif_2_land_1_lpi_1_dfm;
  reg aif_3_land_lpi_1_dfm;
  reg if_5_if_nbw_stat_sva;
  reg else_8_land_lpi_1_dfm;
  reg I_write_flag_sva;
  reg W_write_flag_sva;
  reg [1:0] skid_buf_top_cnt_sva_1_1;
  wire [2:0] nl_skid_buf_top_cnt_sva_1_1;
  reg [15:0] mac_data_data_sva_dfm_2_1;
  reg [4:0] I_vld_pntr_sva_dfm_1_1;
  reg [4:0] W_vld_pntr_sva_dfm_1_1;
  wire O_rd_data_rsci_idat_mx0c0;
  wire O_rd_data_rsci_idat_mx0c1;
  wire O_rd_data_rsci_idat_mx0c2;
  wire [15:0] O_write_data_data_sva_mx0;
  wire skid_buf_top_wr_ptr_sva_0_mx0w0;
  wire skid_buf_top_wr_ptr_sva_1_mx0w0;
  wire [49:0] O_instr_in_crt_lpi_1_dfm_mx0;
  wire O_data_vld_sva_mx0c1;
  wire else_8_land_lpi_1_dfm_mx0w0;
  wire [15:0] mac_data_data_sva_dfm_3;
  wire skid_buf_top_push_and_psp_1;
  wire [49:0] I_instr_in_crt_lpi_1_dfm_1_mx0;
  wire [49:0] W_instr_in_crt_lpi_1_dfm_1_mx0;
  wire flags_top_1_1_sva_mx0c1;
  wire skid_buf_top_push_nor_psp_mx0w0;
  wire skid_buf_top_push_and_1_psp_mx0w0;
  wire [4:0] O_mac_tile_bound_4_lpi_1_dfm_mx0;
  wire [4:0] O_mac_tile_bound_3_lpi_1_dfm_mx0;
  wire [4:0] O_mac_tile_bound_2_lpi_1_dfm_mx0;
  wire [4:0] O_mac_tile_bound_1_lpi_1_dfm_mx0;
  wire [4:0] O_mac_tile_bound_0_lpi_1_dfm_mx0;
  wire [4:0] O_vld_zg_pntr_sva_4;
  wire [5:0] nl_O_vld_zg_pntr_sva_4;
  wire skid_buf_top_peek_nor_m1c_1;
  wire skid_buf_top_peek_and_m1c_2;
  wire skid_buf_top_peek_and_m1c_3;
  wire O_data_vld_sva_dfm_4_mx0w0;
  wire if_5_and_1_m1c_1;
  wire if_5_if_5_nor_m1c_1;
  wire [4:0] I_wr_pntr_sva_dfm_1;
  wire [4:0] W_wr_pntr_sva_dfm_1;
  wire [1:0] skid_buf_wr_zero_guard_cnt_sva_5;
  wire [2:0] nl_skid_buf_wr_zero_guard_cnt_sva_5;
  wire [4:0] W_mac_tile_bound_4_lpi_1_dfm_mx0;
  wire [4:0] W_mac_tile_bound_3_lpi_1_dfm_mx0;
  wire [4:0] W_mac_tile_bound_2_lpi_1_dfm_mx0;
  wire [4:0] W_mac_tile_bound_1_lpi_1_dfm_mx0;
  wire [4:0] W_mac_tile_bound_0_lpi_1_dfm_mx0;
  wire [4:0] I_mac_tile_bound_4_lpi_1_dfm_mx0;
  wire [4:0] I_mac_tile_bound_3_lpi_1_dfm_mx0;
  wire [4:0] I_mac_tile_bound_2_lpi_1_dfm_mx0;
  wire [4:0] I_mac_tile_bound_1_lpi_1_dfm_mx0;
  wire [4:0] I_mac_tile_bound_0_lpi_1_dfm_mx0;
  wire [4:0] libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_18;
  wire libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_21;
  wire libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_22;
  wire libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_23;
  wire [24:0] libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_24;
  wire [24:0] libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_25;
  wire [4:0] libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_19;
  wire libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_26;
  wire libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_27;
  wire libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_28;
  wire [24:0] libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_29;
  wire [24:0] libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_30;
  wire [4:0] libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_20;
  wire libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_31;
  wire libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_32;
  wire libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_33;
  wire [24:0] libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_34;
  wire [24:0] libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_35;
  reg reg_W_instr_in_rsci_oswt_cse_1;
  wire skid_buf_top_cnt_and_1_cse;
  wire nand_73_cse;
  wire and_331_cse;
  wire and_dcpl_34;
  wire or_dcpl;
  wire [1:0] skid_buf_top_push_1_acc_1_tmp;
  wire [2:0] nl_skid_buf_top_push_1_acc_1_tmp;
  wire or_tmp_299;
  wire or_tmp_300;
  wire not_tmp_156;
  wire nand_tmp;
  wire mux_tmp_245;
  wire mux_tmp_247;
  wire mux_tmp_251;
  wire not_tmp_165;
  wire nand_tmp_39;
  wire not_tmp_172;
  wire nand_tmp_46;
  wire and_dcpl_58;
  wire nor_tmp_182;
  wire and_tmp_102;
  wire and_tmp_103;
  wire and_tmp_104;
  wire nor_tmp_189;
  wire and_tmp_107;
  wire mux_tmp_296;
  wire not_tmp_191;
  wire not_tmp_193;
  wire nor_tmp_217;
  wire mux_404_tmp;
  wire and_370_cse;
  wire and_541_cse;
  wire nand_129_cse;
  wire and_526_cse;
  wire and_432_cse;
  wire and_544_cse;
  wire nor_215_cse;
  wire or_756_cse;
  wire or_601_cse;
  wire or_600_cse;
  wire or_598_cse;
  wire nor_303_cse;
  wire or_620_cse;
  wire and_395_cse;
  wire and_426_cse;
  wire skid_buf_top_pop_skid_buf_top_pop_and_4_itm;
  wire skid_buf_top_pop_skid_buf_top_pop_and_2_itm;
  wire mux_530_itm;
  wire mux_543_itm;
  wire mux_642_itm;
  wire mux_663_itm;
  wire skid_buf_top_rd_ptr_and_cse;

  wire[0:0] mux_355_nl;
  wire[0:0] mux_354_nl;
  wire[0:0] nor_182_nl;
  wire[0:0] nor_183_nl;
  wire[0:0] mux_353_nl;
  wire[0:0] nor_184_nl;
  wire[0:0] nor_185_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] nor_178_nl;
  wire[0:0] nor_179_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] nor_180_nl;
  wire[0:0] nor_181_nl;
  wire[0:0] if_5_if_or_nl;
  wire[0:0] if_5_if_or_2_nl;
  wire[0:0] if_5_if_or_3_nl;
  wire[0:0] if_5_if_or_4_nl;
  wire[0:0] if_5_if_or_5_nl;
  wire[0:0] mux_388_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] mux_386_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] or_97_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] and_293_nl;
  wire[0:0] and_294_nl;
  wire[0:0] mux_419_nl;
  wire[0:0] nor_175_nl;
  wire[0:0] mux_418_nl;
  wire[0:0] nand_37_nl;
  wire[0:0] nand_36_nl;
  wire[0:0] mux_428_nl;
  wire[0:0] and_302_nl;
  wire[0:0] mux_430_nl;
  wire[0:0] and_301_nl;
  wire[0:0] mux_432_nl;
  wire[0:0] and_300_nl;
  wire[0:0] mux_597_nl;
  wire[0:0] mux_596_nl;
  wire[0:0] mux_595_nl;
  wire[0:0] or_593_nl;
  wire[0:0] mux_601_nl;
  wire[0:0] and_537_nl;
  wire[0:0] nor_302_nl;
  wire[0:0] mux_600_nl;
  wire[0:0] mux_599_nl;
  wire[0:0] nand_101_nl;
  wire[0:0] nand_100_nl;
  wire[0:0] mux_605_nl;
  wire[0:0] and_533_nl;
  wire[0:0] nor_299_nl;
  wire[0:0] mux_604_nl;
  wire[0:0] mux_603_nl;
  wire[0:0] nand_108_nl;
  wire[0:0] nand_107_nl;
  wire[0:0] mux_614_nl;
  wire[0:0] mux_613_nl;
  wire[0:0] and_388_nl;
  wire[0:0] and_387_nl;
  wire[0:0] mux_612_nl;
  wire[0:0] mux_611_nl;
  wire[0:0] mux_610_nl;
  wire[0:0] mux_609_nl;
  wire[0:0] and_385_nl;
  wire[0:0] and_384_nl;
  wire[0:0] mux_608_nl;
  wire[0:0] mux_607_nl;
  wire[0:0] mux_606_nl;
  wire[0:0] mux_459_nl;
  wire[0:0] mux_458_nl;
  wire[0:0] mux_457_nl;
  wire[0:0] mux_456_nl;
  wire[0:0] else_8_else_8_or_2_nl;
  wire[0:0] mux_490_nl;
  wire[0:0] mux_489_nl;
  wire[0:0] mux_488_nl;
  wire[0:0] mux_487_nl;
  wire[0:0] mux_517_nl;
  wire[0:0] mux_516_nl;
  wire[0:0] mux_515_nl;
  wire[0:0] mux_514_nl;
  wire[0:0] mux_618_nl;
  wire[0:0] and_393_nl;
  wire[0:0] mux_617_nl;
  wire[0:0] and_392_nl;
  wire[0:0] if_6_if_6_and_3_nl;
  wire[0:0] if_6_if_6_and_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] mux_340_nl;
  wire[0:0] and_52_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] and_49_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] if_6_if_6_and_9_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] mux_646_nl;
  wire[0:0] mux_645_nl;
  wire[0:0] mux_719_nl;
  wire[0:0] mux_644_nl;
  wire[0:0] mux_720_nl;
  wire[0:0] mux_643_nl;
  wire[0:0] or_531_nl;
  wire[0:0] mux_553_nl;
  wire[0:0] or_555_nl;
  wire[0:0] or_556_nl;
  wire[0:0] mux_672_nl;
  wire[0:0] mux_671_nl;
  wire[0:0] mux_670_nl;
  wire[0:0] mux_716_nl;
  wire[0:0] mux_669_nl;
  wire[0:0] mux_668_nl;
  wire[0:0] mux_667_nl;
  wire[0:0] mux_666_nl;
  wire[0:0] mux_721_nl;
  wire[0:0] mux_665_nl;
  wire[0:0] mux_722_nl;
  wire[0:0] mux_664_nl;
  wire[0:0] mux_675_nl;
  wire[0:0] or_757_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] if_6_mux_3_nl;
  wire[0:0] if_6_if_if_6_if_and_nl;
  wire[0:0] mux_561_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] and_172_nl;
  wire[0:0] mux_558_nl;
  wire[0:0] and_169_nl;
  wire[0:0] mux_556_nl;
  wire[0:0] mux_555_nl;
  wire[0:0] mux_717_nl;
  wire[0:0] mux_718_nl;
  wire[0:0] skid_buf_top_push_1_skid_buf_top_push_1_and_nl;
  wire[0:0] skid_buf_top_push_1_skid_buf_top_push_1_and_1_nl;
  wire[0:0] nand_85_nl;
  wire[15:0] UPDATE_PSUM_acc_nl;
  wire[16:0] nl_UPDATE_PSUM_acc_nl;
  wire[15:0] UPDATE_PSUM_mux_8_nl;
  wire[15:0] UPDATE_PSUM_mux_9_nl;
  wire[0:0] and_550_nl;
  wire[0:0] and_3_nl;
  wire[0:0] else_3_aelse_mux_1_nl;
  wire[0:0] and_125_nl;
  wire[0:0] aelse_2_aelse_2_and_2_nl;
  wire[0:0] aelse_3_aelse_3_and_nl;
  wire[1:0] skid_buf_wr_zero_guard_pop_acc_nl;
  wire[2:0] nl_skid_buf_wr_zero_guard_pop_acc_nl;
  wire[0:0] nor_nl;
  wire[0:0] mux_562_nl;
  wire[0:0] mux_563_nl;
  wire[4:0] if_if_mux_1_nl;
  wire[0:0] if_6_if_if_not_5_nl;
  wire[0:0] if_6_mux_4_nl;
  wire[0:0] if_6_else_mux_2_nl;
  wire[0:0] if_6_else_if_if_6_else_if_or_nl;
  wire[0:0] if_7_mux_3_nl;
  wire[0:0] if_7_mux_1_nl;
  wire[4:0] O_mac_pntr_mux_1_nl;
  wire[4:0] O_vld_zg_pntr_mux_1_nl;
  wire[0:0] O_vld_zg_pntr_and_nl;
  wire[4:0] mux_5_nl;
  wire[0:0] asn_I_wr_pntr_sva_nand_nl;
  wire[4:0] mux_3_nl;
  wire[0:0] nand_91_nl;
  wire[0:0] nand_nl;
  wire[0:0] or_590_nl;
  wire[0:0] if_5_and_5_nl;
  wire[0:0] if_5_and_4_nl;
  wire[0:0] and_51_nl;
  wire[0:0] and_50_nl;
  wire[0:0] and_54_nl;
  wire[0:0] and_53_nl;
  wire[0:0] and_58_nl;
  wire[0:0] and_56_nl;
  wire[0:0] mux_345_nl;
  wire[0:0] nand_83_nl;
  wire[0:0] nand_84_nl;
  wire[0:0] and_64_nl;
  wire[0:0] and_63_nl;
  wire[0:0] mux_356_nl;
  wire[0:0] and_75_nl;
  wire[0:0] and_74_nl;
  wire[0:0] and_92_nl;
  wire[0:0] and_91_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] mux_368_nl;
  wire[0:0] nand_14_nl;
  wire[0:0] nand_13_nl;
  wire[0:0] and_305_nl;
  wire[0:0] nor_208_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] nor_203_nl;
  wire[0:0] nor_204_nl;
  wire[0:0] mux_397_nl;
  wire[0:0] or_119_nl;
  wire[0:0] or_117_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] mux_402_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] nand_75_nl;
  wire[0:0] or_192_nl;
  wire[0:0] or_191_nl;
  wire[0:0] nand_31_nl;
  wire[0:0] nand_32_nl;
  wire[0:0] nand_34_nl;
  wire[0:0] nand_33_nl;
  wire[0:0] mux_414_nl;
  wire[0:0] mux_413_nl;
  wire[0:0] nand_35_nl;
  wire[0:0] mux_416_nl;
  wire[0:0] mux_415_nl;
  wire[0:0] and_128_nl;
  wire[0:0] and_127_nl;
  wire[0:0] mux_425_nl;
  wire[0:0] and_129_nl;
  wire[0:0] mux_423_nl;
  wire[0:0] and_126_nl;
  wire[0:0] or_267_nl;
  wire[0:0] mux_421_nl;
  wire[0:0] nor_201_nl;
  wire[0:0] nor_200_nl;
  wire[0:0] nor_199_nl;
  wire[0:0] mux_445_nl;
  wire[0:0] nor_195_nl;
  wire[0:0] nor_196_nl;
  wire[0:0] mux_443_nl;
  wire[0:0] or_394_nl;
  wire[0:0] or_392_nl;
  wire[0:0] mux_461_nl;
  wire[0:0] or_422_nl;
  wire[0:0] or_421_nl;
  wire[0:0] mux_465_nl;
  wire[0:0] mux_464_nl;
  wire[0:0] mux_463_nl;
  wire[0:0] nor_191_nl;
  wire[0:0] nor_192_nl;
  wire[0:0] mux_466_nl;
  wire[0:0] and_299_nl;
  wire[0:0] mux_475_nl;
  wire[0:0] mux_474_nl;
  wire[0:0] or_428_nl;
  wire[0:0] mux_473_nl;
  wire[0:0] mux_472_nl;
  wire[0:0] mux_471_nl;
  wire[0:0] mux_470_nl;
  wire[0:0] mux_469_nl;
  wire[0:0] mux_468_nl;
  wire[0:0] or_425_nl;
  wire[0:0] mux_485_nl;
  wire[0:0] mux_484_nl;
  wire[0:0] or_434_nl;
  wire[0:0] mux_483_nl;
  wire[0:0] mux_482_nl;
  wire[0:0] mux_481_nl;
  wire[0:0] mux_480_nl;
  wire[0:0] mux_479_nl;
  wire[0:0] mux_478_nl;
  wire[0:0] or_431_nl;
  wire[0:0] mux_493_nl;
  wire[0:0] nor_190_nl;
  wire[0:0] mux_502_nl;
  wire[0:0] mux_501_nl;
  wire[0:0] or_445_nl;
  wire[0:0] mux_500_nl;
  wire[0:0] mux_499_nl;
  wire[0:0] mux_498_nl;
  wire[0:0] mux_497_nl;
  wire[0:0] mux_496_nl;
  wire[0:0] mux_495_nl;
  wire[0:0] or_442_nl;
  wire[0:0] mux_512_nl;
  wire[0:0] mux_511_nl;
  wire[0:0] or_451_nl;
  wire[0:0] mux_510_nl;
  wire[0:0] mux_509_nl;
  wire[0:0] mux_508_nl;
  wire[0:0] mux_507_nl;
  wire[0:0] mux_506_nl;
  wire[0:0] mux_505_nl;
  wire[0:0] or_448_nl;
  wire[0:0] and_153_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] mux_519_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] mux_534_nl;
  wire[0:0] mux_533_nl;
  wire[0:0] mux_532_nl;
  wire[0:0] mux_531_nl;
  wire[0:0] and_171_nl;
  wire[0:0] and_170_nl;
  wire[0:0] and_296_nl;
  wire[0:0] and_297_nl;
  wire[0:0] mux_570_nl;
  wire[0:0] mux_569_nl;
  wire[0:0] and_175_nl;
  wire[0:0] and_174_nl;
  wire[0:0] mux_568_nl;
  wire[0:0] mux_567_nl;
  wire[0:0] mux_566_nl;
  wire[0:0] or_493_nl;
  wire[0:0] mux_572_nl;
  wire[0:0] nor_188_nl;
  wire[0:0] nor_189_nl;
  wire[0:0] mux_374_nl;
  wire[0:0] mux_373_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] mux_371_nl;
  wire[0:0] and_95_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] nand_16_nl;
  wire[0:0] mux_381_nl;
  wire[0:0] nand_57_nl;
  wire[0:0] nand_58_nl;
  wire[0:0] mux_529_nl;
  wire[0:0] mux_528_nl;
  wire[0:0] mux_527_nl;
  wire[0:0] nor_138_nl;
  wire[0:0] mux_526_nl;
  wire[0:0] nor_136_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] nor_134_nl;
  wire[0:0] mux_523_nl;
  wire[0:0] nor_130_nl;
  wire[0:0] mux_542_nl;
  wire[0:0] mux_541_nl;
  wire[0:0] mux_540_nl;
  wire[0:0] nor_149_nl;
  wire[0:0] mux_539_nl;
  wire[0:0] nor_147_nl;
  wire[0:0] mux_538_nl;
  wire[0:0] mux_537_nl;
  wire[0:0] nor_145_nl;
  wire[0:0] mux_536_nl;
  wire[0:0] nor_140_nl;
  wire[0:0] mux_585_nl;
  wire[0:0] mux_587_nl;
  wire[0:0] nor_307_nl;
  wire[0:0] and_365_nl;
  wire[0:0] mux_586_nl;
  wire[0:0] nand_96_nl;
  wire[0:0] mux_589_nl;
  wire[0:0] mux_593_nl;
  wire[0:0] mux_592_nl;
  wire[0:0] mux_591_nl;
  wire[0:0] and_539_nl;
  wire[0:0] nor_304_nl;
  wire[0:0] and_535_nl;
  wire[0:0] nor_301_nl;
  wire[0:0] mux_638_nl;
  wire[0:0] mux_637_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] mux_635_nl;
  wire[0:0] mux_641_nl;
  wire[0:0] and_516_nl;
  wire[0:0] and_425_nl;
  wire[0:0] mux_640_nl;
  wire[0:0] mux_662_nl;
  wire[0:0] mux_661_nl;
  wire[15:0] mux_723_nl;
  wire[15:0] UPDATE_PSUM_FROM_TOP_mux_5_nl;
  wire[0:0] UPDATE_PSUM_FROM_TOP_or_2_nl;
  wire[15:0] if_10_mux_97_nl;
  wire[15:0] if_10_mux_98_nl;
  wire[15:0] if_10_mux_99_nl;
  wire[15:0] if_10_mux_100_nl;
  wire[15:0] if_10_mux_101_nl;
  wire[15:0] if_10_mux_102_nl;
  wire[15:0] if_10_mux_103_nl;
  wire[15:0] if_10_mux_104_nl;
  wire[15:0] if_10_mux_105_nl;
  wire[15:0] if_10_mux_106_nl;
  wire[15:0] if_10_mux_107_nl;
  wire[15:0] if_10_mux_108_nl;
  wire[15:0] if_10_mux_109_nl;
  wire[15:0] if_10_mux_110_nl;
  wire[15:0] if_10_mux_111_nl;
  wire[15:0] if_10_mux_112_nl;
  wire[15:0] if_10_mux_113_nl;
  wire[15:0] if_10_mux_114_nl;
  wire[15:0] if_10_mux_115_nl;
  wire[15:0] if_10_mux_116_nl;
  wire[15:0] if_10_mux_117_nl;
  wire[15:0] if_10_mux_118_nl;
  wire[15:0] if_10_mux_119_nl;
  wire[15:0] if_10_mux_120_nl;
  wire[15:0] if_10_mux_121_nl;
  wire[15:0] if_10_mux_122_nl;
  wire[15:0] if_10_mux_123_nl;
  wire[15:0] if_10_mux_124_nl;
  wire[15:0] if_10_mux_125_nl;
  wire[15:0] if_10_mux_126_nl;
  wire[15:0] if_10_mux_127_nl;
  wire[15:0] mux_724_nl;
  wire[15:0] UPDATE_PSUM_FROM_TOP_mux_6_nl;
  wire[0:0] UPDATE_PSUM_FROM_TOP_or_3_nl;
  wire[15:0] if_9_mux_97_nl;
  wire[15:0] if_9_mux_98_nl;
  wire[15:0] if_9_mux_99_nl;
  wire[15:0] if_9_mux_100_nl;
  wire[15:0] if_9_mux_101_nl;
  wire[15:0] if_9_mux_102_nl;
  wire[15:0] if_9_mux_103_nl;
  wire[15:0] if_9_mux_104_nl;
  wire[15:0] if_9_mux_105_nl;
  wire[15:0] if_9_mux_106_nl;
  wire[15:0] if_9_mux_107_nl;
  wire[15:0] if_9_mux_108_nl;
  wire[15:0] if_9_mux_109_nl;
  wire[15:0] if_9_mux_110_nl;
  wire[15:0] if_9_mux_111_nl;
  wire[15:0] if_9_mux_112_nl;
  wire[15:0] if_9_mux_113_nl;
  wire[15:0] if_9_mux_114_nl;
  wire[15:0] if_9_mux_115_nl;
  wire[15:0] if_9_mux_116_nl;
  wire[15:0] if_9_mux_117_nl;
  wire[15:0] if_9_mux_118_nl;
  wire[15:0] if_9_mux_119_nl;
  wire[15:0] if_9_mux_120_nl;
  wire[15:0] if_9_mux_121_nl;
  wire[15:0] if_9_mux_122_nl;
  wire[15:0] if_9_mux_123_nl;
  wire[15:0] if_9_mux_124_nl;
  wire[15:0] if_9_mux_125_nl;
  wire[15:0] if_9_mux_126_nl;
  wire[15:0] if_9_mux_127_nl;
  wire[1:0] skid_buf_top_pop_1_mux_1_nl;
  wire[0:0] and_549_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [24:0] nl_O_mac_pntr_cntInst_run_rg_loop_bound;
  assign nl_O_mac_pntr_cntInst_run_rg_loop_bound = O_instr_in_crt_lpi_1_dfm_mx0[24:0];
  wire [24:0] nl_O_mac_pntr_cntInst_run_rg_tile_sizes;
  assign nl_O_mac_pntr_cntInst_run_rg_tile_sizes = O_instr_in_crt_lpi_1_dfm_mx0[49:25];
  wire [24:0] nl_O_mac_pntr_cntInst_run_rg_counter_in;
  assign nl_O_mac_pntr_cntInst_run_rg_counter_in = {O_mac_counter_4_sva , O_mac_counter_3_sva
      , O_mac_counter_2_sva , O_mac_counter_1_sva , O_mac_counter_0_sva};
  wire [24:0] nl_O_mac_pntr_cntInst_run_rg_tile_bound_in;
  assign nl_O_mac_pntr_cntInst_run_rg_tile_bound_in = {O_mac_tile_bound_4_lpi_1_dfm_mx0
      , O_mac_tile_bound_3_lpi_1_dfm_mx0 , O_mac_tile_bound_2_lpi_1_dfm_mx0 , O_mac_tile_bound_1_lpi_1_dfm_mx0
      , O_mac_tile_bound_0_lpi_1_dfm_mx0};
  wire [24:0] nl_W_mac_pntr_cntInst_run_rg_loop_bound;
  assign nl_W_mac_pntr_cntInst_run_rg_loop_bound = W_instr_in_crt_lpi_1_dfm_1_mx0[24:0];
  wire [24:0] nl_W_mac_pntr_cntInst_run_rg_tile_sizes;
  assign nl_W_mac_pntr_cntInst_run_rg_tile_sizes = W_instr_in_crt_lpi_1_dfm_1_mx0[49:25];
  wire [24:0] nl_W_mac_pntr_cntInst_run_rg_counter_in;
  assign nl_W_mac_pntr_cntInst_run_rg_counter_in = {W_mac_counter_4_sva , W_mac_counter_3_sva
      , W_mac_counter_2_sva , W_mac_counter_1_sva , W_mac_counter_0_sva};
  wire [24:0] nl_W_mac_pntr_cntInst_run_rg_tile_bound_in;
  assign nl_W_mac_pntr_cntInst_run_rg_tile_bound_in = {W_mac_tile_bound_4_lpi_1_dfm_mx0
      , W_mac_tile_bound_3_lpi_1_dfm_mx0 , W_mac_tile_bound_2_lpi_1_dfm_mx0 , W_mac_tile_bound_1_lpi_1_dfm_mx0
      , W_mac_tile_bound_0_lpi_1_dfm_mx0};
  wire [24:0] nl_I_mac_pntr_cntInst_run_rg_loop_bound;
  assign nl_I_mac_pntr_cntInst_run_rg_loop_bound = I_instr_in_crt_lpi_1_dfm_1_mx0[24:0];
  wire [24:0] nl_I_mac_pntr_cntInst_run_rg_tile_sizes;
  assign nl_I_mac_pntr_cntInst_run_rg_tile_sizes = I_instr_in_crt_lpi_1_dfm_1_mx0[49:25];
  wire [24:0] nl_I_mac_pntr_cntInst_run_rg_counter_in;
  assign nl_I_mac_pntr_cntInst_run_rg_counter_in = {I_mac_counter_4_sva , I_mac_counter_3_sva
      , I_mac_counter_2_sva , I_mac_counter_1_sva , I_mac_counter_0_sva};
  wire [24:0] nl_I_mac_pntr_cntInst_run_rg_tile_bound_in;
  assign nl_I_mac_pntr_cntInst_run_rg_tile_bound_in = {I_mac_tile_bound_4_lpi_1_dfm_mx0
      , I_mac_tile_bound_3_lpi_1_dfm_mx0 , I_mac_tile_bound_2_lpi_1_dfm_mx0 , I_mac_tile_bound_1_lpi_1_dfm_mx0
      , I_mac_tile_bound_0_lpi_1_dfm_mx0};
  O_addr_cnt_5_O_addr_type_L1_1  O_mac_pntr_cntInst_run_rg (
      .loop_bound(nl_O_mac_pntr_cntInst_run_rg_loop_bound[24:0]),
      .tile_sizes(nl_O_mac_pntr_cntInst_run_rg_tile_sizes[24:0]),
      .pntr_in(O_mac_pntr_sva),
      .pntr_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_18),
      .irrel_at_max_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_21),
      .irrel_at_zero_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_22),
      .all_at_max_1_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_23),
      .counter_in(nl_O_mac_pntr_cntInst_run_rg_counter_in[24:0]),
      .counter_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_24),
      .tile_bound_in(nl_O_mac_pntr_cntInst_run_rg_tile_bound_in[24:0]),
      .tile_bound_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_25)
    );
  O_addr_cnt_5_O_addr_type_L1_1  W_mac_pntr_cntInst_run_rg (
      .loop_bound(nl_W_mac_pntr_cntInst_run_rg_loop_bound[24:0]),
      .tile_sizes(nl_W_mac_pntr_cntInst_run_rg_tile_sizes[24:0]),
      .pntr_in(W_mac_pntr_sva),
      .pntr_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_19),
      .irrel_at_max_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_26),
      .irrel_at_zero_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_27),
      .all_at_max_1_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_28),
      .counter_in(nl_W_mac_pntr_cntInst_run_rg_counter_in[24:0]),
      .counter_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_29),
      .tile_bound_in(nl_W_mac_pntr_cntInst_run_rg_tile_bound_in[24:0]),
      .tile_bound_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_30)
    );
  O_addr_cnt_5_O_addr_type_L1_1  I_mac_pntr_cntInst_run_rg (
      .loop_bound(nl_I_mac_pntr_cntInst_run_rg_loop_bound[24:0]),
      .tile_sizes(nl_I_mac_pntr_cntInst_run_rg_tile_sizes[24:0]),
      .pntr_in(I_mac_pntr_sva),
      .pntr_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_20),
      .irrel_at_max_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_31),
      .irrel_at_zero_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_32),
      .all_at_max_1_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_33),
      .counter_in(nl_I_mac_pntr_cntInst_run_rg_counter_in[24:0]),
      .counter_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_34),
      .tile_bound_in(nl_I_mac_pntr_cntInst_run_rg_tile_bound_in[24:0]),
      .tile_bound_out(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_35)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_wr_data_rsci
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_wr_data_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .O_wr_data_rsc_dat(O_wr_data_rsc_dat),
      .O_wr_data_rsc_vld(O_wr_data_rsc_vld),
      .O_wr_data_rsc_rdy(O_wr_data_rsc_rdy),
      .run_wen(run_wen),
      .O_wr_data_rsci_oswt(reg_O_wr_data_rsci_irdy_run_psct_cse),
      .run_wten(run_wten),
      .O_wr_data_rsci_ivld_mxwt(O_wr_data_rsci_ivld_mxwt),
      .O_wr_data_rsci_idat_mxwt(O_wr_data_rsci_idat_mxwt)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_rd_data_rsci
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_rd_data_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .O_rd_data_rsc_dat(O_rd_data_rsc_dat),
      .O_rd_data_rsc_vld(O_rd_data_rsc_vld),
      .O_rd_data_rsc_rdy(O_rd_data_rsc_rdy),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .O_rd_data_rsci_oswt(reg_O_rd_data_rsci_ivld_run_psct_cse),
      .O_rd_data_rsci_irdy_mxwt(O_rd_data_rsci_irdy_mxwt),
      .O_rd_data_rsci_idat(O_rd_data_rsci_idat)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_wr_data_rsci
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_wr_data_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .I_wr_data_rsc_dat(I_wr_data_rsc_dat),
      .I_wr_data_rsc_vld(I_wr_data_rsc_vld),
      .I_wr_data_rsc_rdy(I_wr_data_rsc_rdy),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .I_wr_data_rsci_oswt(reg_I_wr_data_rsci_irdy_run_psct_cse),
      .I_wr_data_rsci_ivld_mxwt(I_wr_data_rsci_ivld_mxwt),
      .I_wr_data_rsci_idat_mxwt(I_wr_data_rsci_idat_mxwt)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_wr_data_rsci
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_wr_data_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .W_wr_data_rsc_dat(W_wr_data_rsc_dat),
      .W_wr_data_rsc_vld(W_wr_data_rsc_vld),
      .W_wr_data_rsc_rdy(W_wr_data_rsc_rdy),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .W_wr_data_rsci_oswt(reg_W_wr_data_rsci_irdy_run_psct_cse),
      .W_wr_data_rsci_ivld_mxwt(W_wr_data_rsci_ivld_mxwt),
      .W_wr_data_rsci_idat_mxwt(W_wr_data_rsci_idat_mxwt)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_wr_data_zero_guard_rsci
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_wr_data_zero_guard_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .wr_data_zero_guard_rsc_dat(wr_data_zero_guard_rsc_dat),
      .wr_data_zero_guard_rsc_vld(wr_data_zero_guard_rsc_vld),
      .wr_data_zero_guard_rsc_rdy(wr_data_zero_guard_rsc_rdy),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .wr_data_zero_guard_rsci_oswt(reg_wr_data_zero_guard_rsci_oswt_cse),
      .wr_data_zero_guard_rsci_ivld_mxwt(wr_data_zero_guard_rsci_ivld_mxwt),
      .wr_data_zero_guard_rsci_idat_mxwt(wr_data_zero_guard_rsci_idat_mxwt)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_instr_in_rsci
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_O_instr_in_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .O_instr_in_rsc_dat(O_instr_in_rsc_dat),
      .O_instr_in_rsc_vld(O_instr_in_rsc_vld),
      .O_instr_in_rsc_rdy(O_instr_in_rsc_rdy),
      .run_wen(run_wen),
      .O_instr_in_rsci_oswt(reg_W_instr_in_rsci_oswt_cse_1),
      .O_instr_in_rsci_wen_comp(O_instr_in_rsci_wen_comp),
      .O_instr_in_rsci_idat_mxwt(O_instr_in_rsci_idat_mxwt)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_instr_in_rsci
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_I_instr_in_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .I_instr_in_rsc_dat(I_instr_in_rsc_dat),
      .I_instr_in_rsc_vld(I_instr_in_rsc_vld),
      .I_instr_in_rsc_rdy(I_instr_in_rsc_rdy),
      .run_wen(run_wen),
      .I_instr_in_rsci_oswt(reg_W_instr_in_rsci_oswt_cse_1),
      .I_instr_in_rsci_wen_comp(I_instr_in_rsci_wen_comp),
      .I_instr_in_rsci_idat_mxwt(I_instr_in_rsci_idat_mxwt)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_instr_in_rsci
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_W_instr_in_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .W_instr_in_rsc_dat(W_instr_in_rsc_dat),
      .W_instr_in_rsc_vld(W_instr_in_rsc_vld),
      .W_instr_in_rsc_rdy(W_instr_in_rsc_rdy),
      .run_wen(run_wen),
      .W_instr_in_rsci_oswt(reg_W_instr_in_rsci_oswt_cse_1),
      .W_instr_in_rsci_wen_comp(W_instr_in_rsci_wen_comp),
      .W_instr_in_rsci_idat_mxwt(W_instr_in_rsci_idat_mxwt)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_staller
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .O_instr_in_rsci_wen_comp(O_instr_in_rsci_wen_comp),
      .I_instr_in_rsci_wen_comp(I_instr_in_rsci_wen_comp),
      .W_instr_in_rsci_wen_comp(W_instr_in_rsci_wen_comp)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_run_fsm
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_run_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign or_557_cse = and_295_cse | I_data_vld_sva_dfm_1_1;
  assign flags_wr_zero_guard_and_cse = run_wen & (~ (fsm_output[0]));
  assign operator_2_false_5_operator_2_false_5_operator_2_false_5_or_cse = (mux1h_1_tmp!=2'b00);
  assign W_mac_pntr_and_cse = run_wen & (~(mux_tmp_76 | (fsm_output[0])));
  assign and_302_nl = if_5_and_svs_1 & skid_buf_top_push_nor_psp;
  assign mux_428_nl = MUX_s_1_2_2(mux_tmp_94, and_302_nl, if_5_else_or_tmp_2);
  assign or_359_cse = (~ mux_428_nl) | or_dcpl_226;
  assign and_301_nl = if_5_and_svs_1 & skid_buf_top_push_and_psp;
  assign mux_430_nl = MUX_s_1_2_2(mux_tmp_96, and_301_nl, if_5_else_or_tmp_2);
  assign or_363_cse = (~ mux_430_nl) | or_dcpl_226;
  assign and_300_nl = if_5_and_svs_1 & skid_buf_top_push_and_1_psp;
  assign mux_432_nl = MUX_s_1_2_2(mux_tmp_98, and_300_nl, if_5_else_or_tmp_2);
  assign or_367_cse = (~ mux_432_nl) | or_dcpl_226;
  assign skid_buf_top_rd_ptr_and_cse = or_dcpl & O_rd_data_rsci_irdy_mxwt & and_dcpl_34
      & run_wen & or_570_cse;
  assign and_541_cse = W_wr_data_rsci_ivld_mxwt & if_10_if_equal_1_tmp;
  assign and_370_cse = ((~(operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1_1
      | O_rd_data_rsci_irdy_mxwt)) | if_5_and_svs_1) & and_dcpl_34 & run_wen;
  assign nor_303_cse = ~(and_541_cse | W_data_vld_sva_dfm_1_1 | oif_2_unequal_tmp);
  assign and_526_cse = O_mac_irrel_at_max_sva & flags_top_1_1_sva;
  assign or_620_cse = and_541_cse | W_data_vld_sva_dfm_1_1 | oif_2_unequal_tmp;
  assign mux_459_nl = MUX_s_1_2_2(or_400_cse, or_401_cse, skid_buf_wr_zero_guard_rd_ptr_sva);
  assign mux_457_nl = MUX_s_1_2_2(or_399_cse, or_401_cse, skid_buf_wr_zero_guard_rd_ptr_sva);
  assign mux_456_nl = MUX_s_1_2_2(or_400_cse, or_399_cse, skid_buf_wr_zero_guard_rd_ptr_sva);
  assign mux_458_nl = MUX_s_1_2_2(mux_457_nl, mux_456_nl, skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_460_cse = MUX_s_1_2_2(mux_459_nl, mux_458_nl, nor_tmp_39);
  assign nor_108_cse = ~(land_lpi_1_dfm_1 | (~ if_6_else_if_equal_tmp));
  assign W_mac_irrel_at_maxBuf_and_cse = run_wen & (~((~ reg_W_instr_in_rsci_oswt_cse_1)
      & mux_tmp_76));
  assign nand_129_cse = ~(O_mac_irrel_at_max_sva & flags_top_1_1_sva);
  assign and_393_nl = oif_2_unequal_tmp & or_1_cse & oif_1_unequal_tmp;
  assign and_392_nl = W_wr_data_rsci_ivld_mxwt & if_10_if_equal_1_tmp & mux_343_cse;
  assign mux_617_nl = MUX_s_1_2_2(and_392_nl, mux_343_cse, or_tmp_300);
  assign mux_618_nl = MUX_s_1_2_2(and_393_nl, mux_617_nl, main_stage_0_2);
  assign and_395_cse = ((mux_618_nl & nand_129_cse) | reg_W_instr_in_rsci_oswt_cse_1)
      & run_wen;
  assign skid_buf_top_cnt_and_1_cse = run_wen & and_dcpl;
  assign mux_719_nl = MUX_s_1_2_2(not_tmp_193, mux_642_itm, or_620_cse);
  assign mux_645_nl = MUX_s_1_2_2(not_tmp_193, mux_719_nl, mux_124_itm_1);
  assign mux_720_nl = MUX_s_1_2_2(not_tmp_193, mux_642_itm, or_620_cse);
  assign mux_644_nl = MUX_s_1_2_2(not_tmp_193, mux_720_nl, O_wr_data_rsci_ivld_mxwt);
  assign mux_646_nl = MUX_s_1_2_2(mux_645_nl, mux_644_nl, land_9_lpi_1_dfm_1_1);
  assign mux_643_nl = MUX_s_1_2_2(not_tmp_193, mux_642_itm, or_620_cse);
  assign mux_647_nl = MUX_s_1_2_2(mux_646_nl, mux_643_nl, or_1_cse);
  assign and_426_cse = mux_647_nl & run_wen & main_stage_0_2;
  assign and_544_cse = or_1_cse & oif_1_unequal_tmp;
  assign and_432_cse = wr_data_zero_guard_rsci_ivld_mxwt & (~ flags_wr_zero_guard_sva);
  assign mux_554_cse = MUX_s_1_2_2(or_18_cse, or_tmp_2, main_stage_0_2);
  assign and_172_nl = or_558_cse & mux_tmp_226;
  assign mux_560_nl = MUX_s_1_2_2(and_172_nl, mux_tmp_226, oif_2_unequal_tmp);
  assign and_169_nl = or_558_cse & mux_tmp_224;
  assign mux_555_nl = MUX_s_1_2_2(and_tmp_93, and_tmp, I_data_vld_sva_dfm_1_1);
  assign mux_556_nl = MUX_s_1_2_2(mux_555_nl, mux_554_cse, oif_1_unequal_tmp);
  assign mux_558_nl = MUX_s_1_2_2(and_169_nl, mux_556_nl, oif_2_unequal_tmp);
  assign mux_561_nl = MUX_s_1_2_2(mux_560_nl, mux_558_nl, or_1_cse);
  assign skid_buf_top_push_and_2_cse = run_wen & (~((~ mux_561_nl) | or_dcpl_11 |
      (fsm_output[0])));
  assign or_558_cse = and_541_cse | W_data_vld_sva_dfm_1_1;
  assign and_295_cse = if_9_if_equal_1_tmp & I_wr_data_rsci_ivld_mxwt;
  assign else_3_land_lpi_1_dfm_mx0w0 = land_lpi_1_dfm_1 & land_2_lpi_1_dfm_2;
  assign mux_420_cse = MUX_s_1_2_2(mux_124_itm_1, O_wr_data_rsci_ivld_mxwt, land_9_lpi_1_dfm_1_1);
  assign O_write_data_data_sva_mx0 = MUX_v_16_2_2(O_write_data_data_sva, O_wr_data_rsci_idat_mxwt,
      land_9_lpi_1_dfm_1_1);
  assign or_570_cse = (O_rd_data_rsci_irdy_mxwt & operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1_1
      & and_16_m1c_1) | (if_5_if_nbw_stat_sva_mx1 & and_17_m1c_1);
  assign skid_buf_top_pop_skid_buf_top_pop_and_4_itm = (~ skid_buf_top_rd_ptr_sva_0)
      & skid_buf_top_pop_1_skid_buf_top_pop_1_nand_seb_1;
  assign mux_717_nl = MUX_s_1_2_2(skid_buf_top_rd_ptr_sva_0, skid_buf_top_pop_skid_buf_top_pop_and_4_itm,
      or_570_cse);
  assign skid_buf_top_rd_ptr_sva_0_mx1 = MUX_s_1_2_2(skid_buf_top_rd_ptr_sva_0, mux_717_nl,
      main_stage_0_2);
  assign skid_buf_top_pop_skid_buf_top_pop_and_2_itm = skid_buf_top_pop_1_xor_psp_1
      & skid_buf_top_pop_1_skid_buf_top_pop_1_nand_seb_1;
  assign mux_718_nl = MUX_s_1_2_2(skid_buf_top_rd_ptr_sva_1, skid_buf_top_pop_skid_buf_top_pop_and_2_itm,
      or_570_cse);
  assign skid_buf_top_rd_ptr_sva_1_mx1 = MUX_s_1_2_2(skid_buf_top_rd_ptr_sva_1, mux_718_nl,
      main_stage_0_2);
  assign skid_buf_top_cnt_sva_mx1 = MUX_v_2_2_2(skid_buf_top_cnt_sva, mux1h_7_tmp,
      main_stage_0_2);
  assign skid_buf_top_push_1_skid_buf_top_push_1_and_nl = (~ skid_buf_top_wr_ptr_sva_0)
      & skid_buf_top_push_1_skid_buf_top_push_1_nand_seb_1;
  assign skid_buf_top_wr_ptr_sva_0_mx0w0 = MUX1HOT_s_1_3_2(skid_buf_top_wr_ptr_sva_0,
      skid_buf_top_push_1_skid_buf_top_push_1_and_nl, skid_buf_top_push_nor_psp,
      {nand_11_ssc_1 , and_47_ssc_1 , and_17_m1c_1});
  assign skid_buf_top_wr_ptr_sva_0_mx1 = MUX_s_1_2_2(skid_buf_top_wr_ptr_sva_0, skid_buf_top_wr_ptr_sva_0_mx0w0,
      main_stage_0_2);
  assign skid_buf_top_push_1_skid_buf_top_push_1_and_1_nl = skid_buf_top_push_1_xor_psp_1
      & skid_buf_top_push_1_skid_buf_top_push_1_nand_seb_1;
  assign skid_buf_top_wr_ptr_sva_1_mx0w0 = MUX1HOT_s_1_3_2(skid_buf_top_wr_ptr_sva_1,
      skid_buf_top_push_1_skid_buf_top_push_1_and_1_nl, skid_buf_top_wr_ptr_sva_dfm_1_1,
      {nand_11_ssc_1 , and_47_ssc_1 , and_17_m1c_1});
  assign skid_buf_top_wr_ptr_sva_1_mx1 = MUX_s_1_2_2(skid_buf_top_wr_ptr_sva_1, skid_buf_top_wr_ptr_sva_1_mx0w0,
      main_stage_0_2);
  assign O_instr_in_crt_lpi_1_dfm_mx0 = MUX_v_50_2_2(O_instr_in_crt_lpi_1_dfm, O_instr_in_rsci_idat_mxwt,
      reg_W_instr_in_rsci_oswt_cse_1);
  assign O_write_flag_sva_mx0 = mux_420_cse & main_stage_0_2;
  assign W_data_vld_sva_mx0 = ((if_10_if_equal_1_tmp & W_write_flag_sva_mx0) | W_data_vld_sva_dfm_1_1)
      & main_stage_0_2;
  assign I_data_vld_sva_mx0 = ((if_9_if_equal_1_tmp & I_write_flag_sva_mx0) | I_data_vld_sva_dfm_1_1)
      & main_stage_0_2;
  assign else_8_land_lpi_1_dfm_mx0w0 = land_8_lpi_1_dfm_1 & skid_buf_wr_zero_guard_peek_slc_skid_buf_wr_zero_guard_regs_skid_buf_wr_zero_guard_rd_ptr_1_0_cse_sva_mx0;
  assign else_8_land_lpi_1_dfm_mx1 = MUX_s_1_2_2(else_8_land_lpi_1_dfm_mx0w0, else_8_land_lpi_1_dfm,
      and_dcpl_19);
  assign W_write_flag_sva_mx0 = MUX_s_1_2_2(W_wr_data_rsci_ivld_mxwt, W_write_flag_sva,
      W_data_vld_sva_dfm_1_1);
  assign I_write_flag_sva_mx0 = MUX_s_1_2_2(I_wr_data_rsci_ivld_mxwt, I_write_flag_sva,
      I_data_vld_sva_dfm_1_1);
  assign land_9_lpi_1_dfm_1 = land_8_lpi_1_dfm_1 & (~ skid_buf_wr_zero_guard_peek_slc_skid_buf_wr_zero_guard_regs_skid_buf_wr_zero_guard_rd_ptr_1_0_cse_sva_mx0);
  assign skid_buf_top_pop_1_skid_buf_top_pop_1_nand_seb_1 = ~(skid_buf_top_pop_1_xor_psp_1
      & (~ skid_buf_top_rd_ptr_sva_0));
  assign skid_buf_top_pop_1_xor_psp_1 = skid_buf_top_rd_ptr_sva_0 ^ skid_buf_top_rd_ptr_sva_1;
  assign nand_85_nl = ~(or_svs_1 & if_5_and_svs_1);
  assign if_5_if_nbw_stat_sva_mx1 = MUX_s_1_2_2(O_rd_data_rsci_irdy_mxwt, if_5_if_nbw_stat_sva,
      nand_85_nl);
  assign skid_buf_top_push_1_skid_buf_top_push_1_nand_seb_1 = ~(skid_buf_top_push_1_xor_psp_1
      & (~ skid_buf_top_wr_ptr_sva_0));
  assign skid_buf_top_push_1_xor_psp_1 = skid_buf_top_wr_ptr_sva_0 ^ skid_buf_top_wr_ptr_sva_1;
  assign nand_73_cse = ~(mux_420_cse & main_stage_0_2);
  assign UPDATE_PSUM_mux_9_nl = MUX_v_16_32_2(O_mem_0_sva, O_mem_1_sva, O_mem_2_sva,
      O_mem_3_sva, O_mem_4_sva, O_mem_5_sva, O_mem_6_sva, O_mem_7_sva, O_mem_8_sva,
      O_mem_9_sva, O_mem_10_sva, O_mem_11_sva, O_mem_12_sva, O_mem_13_sva, O_mem_14_sva,
      O_mem_15_sva, O_mem_16_sva, O_mem_17_sva, O_mem_18_sva, O_mem_19_sva, O_mem_20_sva,
      O_mem_21_sva, O_mem_22_sva, O_mem_23_sva, O_mem_24_sva, O_mem_25_sva, O_mem_26_sva,
      O_mem_27_sva, O_mem_28_sva, O_mem_29_sva, O_mem_30_sva, O_mem_31_sva, O_mac_pntr_sva);
  assign and_550_nl = mux_420_cse & main_stage_0_2 & (fsm_output[1]);
  assign UPDATE_PSUM_mux_8_nl = MUX_v_16_2_2(UPDATE_PSUM_mux_9_nl, O_write_data_data_sva_mx0,
      and_550_nl);
  assign nl_UPDATE_PSUM_acc_nl = z_out_2 + UPDATE_PSUM_mux_8_nl;
  assign UPDATE_PSUM_acc_nl = nl_UPDATE_PSUM_acc_nl[15:0];
  assign and_125_nl = nand_73_cse & (~(data_zg_sva & aif_equal_tmp));
  assign else_3_aelse_mux_1_nl = MUX_s_1_2_2(else_3_land_lpi_1_dfm_mx0w0, else_3_land_lpi_1_dfm,
      and_125_nl);
  assign and_3_nl = else_3_aelse_mux_1_nl & (land_lpi_1_dfm_1 | (~ land_2_lpi_1_dfm_2));
  assign mac_data_data_sva_dfm_3 = MUX_v_16_2_2(UPDATE_PSUM_acc_nl, z_out_2, and_3_nl);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1 =
      (skid_buf_top_cnt_sva_mx1!=2'b00);
  assign skid_buf_top_push_and_psp_1 = skid_buf_top_wr_ptr_sva_0_mx1 & (~ skid_buf_top_wr_ptr_sva_1_mx1);
  assign I_instr_in_crt_lpi_1_dfm_1_mx0 = MUX_v_50_2_2(I_instr_in_crt_lpi_1_dfm_1,
      I_instr_in_rsci_idat_mxwt, reg_W_instr_in_rsci_oswt_cse_1);
  assign W_instr_in_crt_lpi_1_dfm_1_mx0 = MUX_v_50_2_2(W_instr_in_crt_lpi_1_dfm_1,
      W_instr_in_rsci_idat_mxwt, reg_W_instr_in_rsci_oswt_cse_1);
  assign or_1_cse = oif_unequal_tmp | O_data_vld_sva;
  assign aelse_2_aelse_2_and_2_nl = lor_2_lpi_1_dfm_1 & lor_1_lpi_1_dfm_1 & or_1_cse;
  assign aif_2_land_1_lpi_1_dfm_mx0 = MUX_s_1_2_2(aelse_2_aelse_2_and_2_nl, aif_2_land_1_lpi_1_dfm,
      and_tmp_56);
  assign aelse_3_aelse_3_and_nl = lor_1_lpi_1_dfm_1 & O_write_flag_sva_mx0;
  assign aif_3_land_lpi_1_dfm_mx0 = MUX_s_1_2_2(aelse_3_aelse_3_and_nl, aif_3_land_lpi_1_dfm,
      and_tmp_56);
  assign mux_124_cse = MUX_v_2_2_2(skid_buf_wr_zero_guard_cnt_sva_5, skid_buf_wr_zero_guard_cnt_sva,
      or_tmp_162);
  assign nl_skid_buf_wr_zero_guard_pop_acc_nl = mux_124_cse + 2'b11;
  assign skid_buf_wr_zero_guard_pop_acc_nl = nl_skid_buf_wr_zero_guard_pop_acc_nl[1:0];
  assign nor_nl = ~(else_8_land_lpi_1_dfm_mx1 | land_9_lpi_1_dfm_1);
  assign mux1h_1_tmp = MUX_v_2_2_2(skid_buf_wr_zero_guard_pop_acc_nl, mux_124_cse,
      nor_nl);
  assign skid_buf_top_push_nor_psp_mx0w0 = ~(skid_buf_top_wr_ptr_sva_0_mx1 | skid_buf_top_wr_ptr_sva_1_mx1);
  assign skid_buf_top_push_and_1_psp_mx0w0 = (~ skid_buf_top_wr_ptr_sva_0_mx1) &
      skid_buf_top_wr_ptr_sva_1_mx1;
  assign nl_if_6_if_3_acc_tmp = ({W_irrel_cnt_sva_4_1 , W_irrel_cnt_sva_0}) + 5'b00001;
  assign if_6_if_3_acc_tmp = nl_if_6_if_3_acc_tmp[4:0];
  assign mux_562_nl = MUX_s_1_2_2(W_mac_irrel_at_maxBuf_sva, if_for_if_for_and_28_tmp,
      reg_W_instr_in_rsci_oswt_cse_1);
  assign W_irrel_cnt_sva_dfm_mx0 = MUX_v_5_2_2(({W_irrel_cnt_sva_4_1 , W_irrel_cnt_sva_0}),
      if_6_if_3_acc_tmp, mux_562_nl);
  assign nl_if_6_if_1_acc_tmp = ({I_irrel_cnt_sva_4_1 , I_irrel_cnt_sva_0}) + 5'b00001;
  assign if_6_if_1_acc_tmp = nl_if_6_if_1_acc_tmp[4:0];
  assign mux_563_nl = MUX_s_1_2_2(I_mac_irrel_at_maxBuf_sva, if_for_if_for_and_27_tmp,
      reg_W_instr_in_rsci_oswt_cse_1);
  assign I_irrel_cnt_sva_dfm_mx0 = MUX_v_5_2_2(({I_irrel_cnt_sva_4_1 , I_irrel_cnt_sva_0}),
      if_6_if_1_acc_tmp, mux_563_nl);
  assign O_mac_tile_bound_4_lpi_1_dfm_mx0 = MUX_v_5_2_2(O_mac_tile_bound_4_lpi_1,
      (O_instr_in_rsci_idat_mxwt[49:45]), reg_W_instr_in_rsci_oswt_cse_1);
  assign O_mac_tile_bound_3_lpi_1_dfm_mx0 = MUX_v_5_2_2(O_mac_tile_bound_3_lpi_1,
      (O_instr_in_rsci_idat_mxwt[44:40]), reg_W_instr_in_rsci_oswt_cse_1);
  assign O_mac_tile_bound_2_lpi_1_dfm_mx0 = MUX_v_5_2_2(O_mac_tile_bound_2_lpi_1,
      (O_instr_in_rsci_idat_mxwt[39:35]), reg_W_instr_in_rsci_oswt_cse_1);
  assign O_mac_tile_bound_1_lpi_1_dfm_mx0 = MUX_v_5_2_2(O_mac_tile_bound_1_lpi_1,
      (O_instr_in_rsci_idat_mxwt[34:30]), reg_W_instr_in_rsci_oswt_cse_1);
  assign O_mac_tile_bound_0_lpi_1_dfm_mx0 = MUX_v_5_2_2(O_mac_tile_bound_0_lpi_1,
      (O_instr_in_rsci_idat_mxwt[29:25]), reg_W_instr_in_rsci_oswt_cse_1);
  assign land_lpi_1_dfm_1 = aif_equal_tmp & data_zg_sva;
  assign nl_O_vld_zg_pntr_sva_4 = O_vld_zg_pntr_sva + 5'b00001;
  assign O_vld_zg_pntr_sva_4 = nl_O_vld_zg_pntr_sva_4[4:0];
  assign if_if_mux_1_nl = MUX_v_5_2_2((O_instr_in_crt_lpi_1_dfm[49:45]), (O_instr_in_rsci_idat_mxwt[49:45]),
      reg_W_instr_in_rsci_oswt_cse_1);
  assign if_6_else_if_equal_tmp = O_vld_zg_pntr_sva_4 == if_if_mux_1_nl;
  assign if_6_if_if_not_5_nl = ~ if_6_else_if_equal_tmp;
  assign if_6_if_if_6_if_and_1_itm = MUX_v_5_2_2(5'b00000, O_vld_zg_pntr_sva_4, if_6_if_if_not_5_nl);
  assign if_6_or_itm = O_write_flag_sva_mx0 | land_lpi_1_dfm_1;
  assign if_6_if_6_mux1h_tmp = MUX_v_5_2_2(O_vld_zg_pntr_sva, if_6_if_if_6_if_and_1_itm,
      if_6_or_itm);
  assign land_2_lpi_1_dfm_2 = (~ O_write_flag_sva_mx0) & aif_2_land_1_lpi_1_dfm_mx0
      & lor_3_lpi_1_dfm_1;
  assign lor_4_lpi_1_dfm_1 = (lor_2_lpi_1_dfm_1 & aif_3_land_lpi_1_dfm_mx0 & lor_3_lpi_1_dfm_1)
      | land_2_lpi_1_dfm_2;
  assign skid_buf_top_peek_nor_m1c_1 = ~(skid_buf_top_rd_ptr_sva_1_mx1 | skid_buf_top_rd_ptr_sva_0_mx1);
  assign skid_buf_top_peek_and_m1c_2 = skid_buf_top_rd_ptr_sva_0_mx1 & (~ skid_buf_top_rd_ptr_sva_1_mx1);
  assign skid_buf_top_peek_and_m1c_3 = skid_buf_top_rd_ptr_sva_1_mx1 & (~ skid_buf_top_rd_ptr_sva_0_mx1);
  assign land_5_lpi_1_dfm_1 = lor_4_lpi_1_dfm_1 & O_mac_irrel_at_max_sva_dfm_mx0;
  assign if_6_else_if_if_6_else_if_or_nl = O_data_vld_sva | if_6_else_if_equal_tmp;
  assign if_6_else_mux_2_nl = MUX_s_1_2_2(O_data_vld_sva, if_6_else_if_if_6_else_if_or_nl,
      O_write_flag_sva_mx0);
  assign if_6_mux_4_nl = MUX_s_1_2_2(if_6_else_mux_2_nl, O_data_vld_sva, land_lpi_1_dfm_1);
  assign O_data_vld_sva_dfm_4_mx0w0 = if_6_mux_4_nl & ((if_6_if_6_mux1h_tmp!=5'b00000)
      | (~(if_6_aif_equal_tmp & libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_21)));
  assign O_data_vld_sva_dfm_4_mx0 = MUX_s_1_2_2(O_data_vld_sva_dfm_4_mx0w0, O_data_vld_sva,
      mux_tmp_76);
  assign if_6_aif_equal_tmp = libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_18
      == if_6_if_6_mux1h_tmp;
  assign if_6_unequal_tmp_2 = ~((W_irrel_cnt_sva_dfm_mx0==5'b00001));
  assign if_6_unequal_tmp_3 = ~((I_irrel_cnt_sva_dfm_mx0==5'b00001));
  assign land_8_lpi_1_dfm_1 = ((mux_124_cse!=2'b00)) & aif_7_equal_tmp & (~ O_data_vld_sva_dfm_4_mx0);
  assign if_7_mux_3_nl = MUX_s_1_2_2(wr_data_zero_guard_rsci_idat_mxwt, skid_buf_wr_zero_guard_regs_0_sva_dfm_1,
      or_dcpl_248);
  assign if_7_mux_1_nl = MUX_s_1_2_2(wr_data_zero_guard_rsci_idat_mxwt, skid_buf_wr_zero_guard_regs_1_sva_dfm_1,
      or_dcpl_246);
  assign skid_buf_wr_zero_guard_peek_slc_skid_buf_wr_zero_guard_regs_skid_buf_wr_zero_guard_rd_ptr_1_0_cse_sva_mx0
      = MUX_s_1_2_2(if_7_mux_3_nl, if_7_mux_1_nl, skid_buf_wr_zero_guard_rd_ptr_sva);
  assign O_mac_pntr_mux_1_nl = MUX_v_5_2_2(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_18,
      O_mac_pntr_sva, and_dcpl_28);
  assign O_vld_zg_pntr_and_nl = if_6_or_itm & (~ and_dcpl_28);
  assign O_vld_zg_pntr_mux_1_nl = MUX_v_5_2_2(O_vld_zg_pntr_sva, if_6_if_if_6_if_and_1_itm,
      O_vld_zg_pntr_and_nl);
  assign aif_7_equal_tmp = O_mac_pntr_mux_1_nl == O_vld_zg_pntr_mux_1_nl;
  assign if_for_if_for_and_28_tmp = (W_instr_in_rsci_idat_mxwt[24:0]==25'b0000100001000010000100001);
  assign if_for_if_for_and_27_tmp = (I_instr_in_rsci_idat_mxwt[24:0]==25'b0000100001000010000100001);
  assign asn_I_wr_pntr_sva_nand_nl = ~(I_wr_data_rsci_ivld_mxwt & main_stage_0_2);
  assign mux_5_nl = MUX_v_5_2_2(I_wr_pntr_sva_dfm_1, I_wr_pntr_sva, asn_I_wr_pntr_sva_nand_nl);
  assign oif_1_unequal_tmp = I_mac_pntr_sva != mux_5_nl;
  assign nand_91_nl = ~(W_wr_data_rsci_ivld_mxwt & main_stage_0_2);
  assign mux_3_nl = MUX_v_5_2_2(W_wr_pntr_sva_dfm_1, W_wr_pntr_sva, nand_91_nl);
  assign oif_2_unequal_tmp = W_mac_pntr_sva != mux_3_nl;
  assign if_5_and_1_m1c_1 = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1_1
      & (~ if_5_and_svs_1);
  assign if_5_if_5_nor_m1c_1 = ~(operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1_1
      | if_5_and_svs_1);
  assign and_17_m1c_1 = if_5_and_svs_1 & or_svs_1;
  assign and_16_m1c_1 = (~ if_5_and_svs_1) & or_svs_1;
  assign nand_11_ssc_1 = ~(or_svs_1 & (~(if_5_else_or_tmp_2 & and_16_m1c_1)));
  assign and_47_ssc_1 = (~ if_5_else_or_tmp_2) & and_16_m1c_1;
  assign if_5_else_or_tmp_2 = O_rd_data_rsci_irdy_mxwt | operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1_1;
  assign I_wr_pntr_sva_dfm_1 = MUX_v_5_2_2(5'b00000, if_9_if_ac_int_cctor_sva_1,
      ((if_9_if_ac_int_cctor_sva_1) != (I_instr_in_crt_lpi_1_dfm_1[49:45])));
  assign if_9_if_equal_1_tmp = I_wr_pntr_sva_dfm_1 == I_vld_pntr_sva_dfm_1_1;
  assign nl_if_9_if_ac_int_cctor_sva_1 = I_wr_pntr_sva + 5'b00001;
  assign if_9_if_ac_int_cctor_sva_1 = nl_if_9_if_ac_int_cctor_sva_1[4:0];
  assign W_wr_pntr_sva_dfm_1 = MUX_v_5_2_2(5'b00000, if_10_if_ac_int_cctor_sva_1,
      ((if_10_if_ac_int_cctor_sva_1) != (W_instr_in_crt_lpi_1_dfm_1[49:45])));
  assign if_10_if_equal_1_tmp = W_wr_pntr_sva_dfm_1 == W_vld_pntr_sva_dfm_1_1;
  assign nl_if_10_if_ac_int_cctor_sva_1 = W_wr_pntr_sva + 5'b00001;
  assign if_10_if_ac_int_cctor_sva_1 = nl_if_10_if_ac_int_cctor_sva_1[4:0];
  assign nl_skid_buf_top_push_1_acc_1_tmp = skid_buf_top_cnt_sva + 2'b01;
  assign skid_buf_top_push_1_acc_1_tmp = nl_skid_buf_top_push_1_acc_1_tmp[1:0];
  assign nand_nl = ~(or_svs_1 & (~(((~ O_rd_data_rsci_irdy_mxwt) & if_5_and_1_m1c_1)
      | (O_rd_data_rsci_irdy_mxwt & if_5_if_5_nor_m1c_1))));
  assign or_590_nl = (O_rd_data_rsci_irdy_mxwt & if_5_and_1_m1c_1 & or_svs_1) | (if_5_if_nbw_stat_sva_mx1
      & if_5_and_svs_1 & or_svs_1);
  assign if_5_and_5_nl = (~ O_rd_data_rsci_irdy_mxwt) & if_5_if_5_nor_m1c_1 & or_svs_1;
  assign if_5_and_4_nl = (~ if_5_if_nbw_stat_sva_mx1) & if_5_and_svs_1 & or_svs_1;
  assign mux1h_7_tmp = MUX1HOT_v_2_4_2(skid_buf_top_cnt_sva, z_out_3, skid_buf_top_push_1_acc_1_tmp,
      skid_buf_top_cnt_sva_1_1, {nand_nl , or_590_nl , if_5_and_5_nl , if_5_and_4_nl});
  assign oif_unequal_tmp = O_mac_pntr_sva != O_vld_zg_pntr_sva;
  assign lor_2_lpi_1_dfm_1 = oif_2_unequal_tmp | W_data_vld_sva_mx0;
  assign lor_1_lpi_1_dfm_1 = oif_1_unequal_tmp | I_data_vld_sva_mx0;
  assign if_for_if_for_and_26_tmp = O_mac_irrel_at_max_sva & (O_instr_in_rsci_idat_mxwt[24:0]==25'b0000100001000010000100001);
  assign O_mac_irrel_at_max_sva_dfm_mx0 = MUX_s_1_2_2(O_mac_irrel_at_max_sva, if_for_if_for_and_26_tmp,
      reg_W_instr_in_rsci_oswt_cse_1);
  assign aif_equal_tmp = O_mac_pntr_sva == O_vld_zg_pntr_sva;
  assign nl_skid_buf_wr_zero_guard_cnt_sva_5 = skid_buf_wr_zero_guard_cnt_sva + 2'b01;
  assign skid_buf_wr_zero_guard_cnt_sva_5 = nl_skid_buf_wr_zero_guard_cnt_sva_5[1:0];
  assign lor_3_lpi_1_dfm_1 = ~(O_mac_irrel_at_max_sva_dfm_mx0 & flags_top_1_1_sva);
  assign W_mac_tile_bound_4_lpi_1_dfm_mx0 = MUX_v_5_2_2(W_mac_tile_bound_4_lpi_1,
      (W_instr_in_rsci_idat_mxwt[49:45]), reg_W_instr_in_rsci_oswt_cse_1);
  assign W_mac_tile_bound_3_lpi_1_dfm_mx0 = MUX_v_5_2_2(W_mac_tile_bound_3_lpi_1,
      (W_instr_in_rsci_idat_mxwt[44:40]), reg_W_instr_in_rsci_oswt_cse_1);
  assign W_mac_tile_bound_2_lpi_1_dfm_mx0 = MUX_v_5_2_2(W_mac_tile_bound_2_lpi_1,
      (W_instr_in_rsci_idat_mxwt[39:35]), reg_W_instr_in_rsci_oswt_cse_1);
  assign W_mac_tile_bound_1_lpi_1_dfm_mx0 = MUX_v_5_2_2(W_mac_tile_bound_1_lpi_1,
      (W_instr_in_rsci_idat_mxwt[34:30]), reg_W_instr_in_rsci_oswt_cse_1);
  assign W_mac_tile_bound_0_lpi_1_dfm_mx0 = MUX_v_5_2_2(W_mac_tile_bound_0_lpi_1,
      (W_instr_in_rsci_idat_mxwt[29:25]), reg_W_instr_in_rsci_oswt_cse_1);
  assign I_mac_tile_bound_4_lpi_1_dfm_mx0 = MUX_v_5_2_2(I_mac_tile_bound_4_lpi_1,
      (I_instr_in_rsci_idat_mxwt[49:45]), reg_W_instr_in_rsci_oswt_cse_1);
  assign I_mac_tile_bound_3_lpi_1_dfm_mx0 = MUX_v_5_2_2(I_mac_tile_bound_3_lpi_1,
      (I_instr_in_rsci_idat_mxwt[44:40]), reg_W_instr_in_rsci_oswt_cse_1);
  assign I_mac_tile_bound_2_lpi_1_dfm_mx0 = MUX_v_5_2_2(I_mac_tile_bound_2_lpi_1,
      (I_instr_in_rsci_idat_mxwt[39:35]), reg_W_instr_in_rsci_oswt_cse_1);
  assign I_mac_tile_bound_1_lpi_1_dfm_mx0 = MUX_v_5_2_2(I_mac_tile_bound_1_lpi_1,
      (I_instr_in_rsci_idat_mxwt[34:30]), reg_W_instr_in_rsci_oswt_cse_1);
  assign I_mac_tile_bound_0_lpi_1_dfm_mx0 = MUX_v_5_2_2(I_mac_tile_bound_0_lpi_1,
      (I_instr_in_rsci_idat_mxwt[29:25]), reg_W_instr_in_rsci_oswt_cse_1);
  assign mux_188_tmp = MUX_v_2_2_2(skid_buf_wr_zero_guard_cnt_sva, skid_buf_wr_zero_guard_cnt_sva_5,
      and_432_cse);
  assign or_tmp_2 = (mux1h_7_tmp!=2'b00);
  assign and_tmp = main_stage_0_2 & or_tmp_2;
  assign and_tmp_1 = if_9_if_equal_1_tmp & I_wr_data_rsci_ivld_mxwt & main_stage_0_2
      & or_tmp_2;
  assign or_tmp_5 = oif_1_unequal_tmp | I_data_vld_sva_dfm_1_1;
  assign mux_tmp_4 = MUX_s_1_2_2(and_tmp_1, and_tmp, or_tmp_5);
  assign and_51_nl = mux_124_itm_1 & mux_tmp_4;
  assign and_50_nl = O_wr_data_rsci_ivld_mxwt & mux_tmp_4;
  assign mux_tmp_6 = MUX_s_1_2_2(and_51_nl, and_50_nl, land_9_lpi_1_dfm_1_1);
  assign or_18_cse = (skid_buf_top_cnt_sva!=2'b00);
  assign or_tmp_10 = and_295_cse | I_data_vld_sva_dfm_1_1 | oif_1_unequal_tmp;
  assign and_54_nl = mux_124_itm_1 & or_tmp_10;
  assign and_53_nl = O_wr_data_rsci_ivld_mxwt & or_tmp_10;
  assign mux_342_cse = MUX_s_1_2_2(and_54_nl, and_53_nl, land_9_lpi_1_dfm_1_1);
  assign mux_343_cse = MUX_s_1_2_2(mux_342_cse, or_tmp_10, or_1_cse);
  assign and_58_nl = oif_2_unequal_tmp & or_1_cse & oif_1_unequal_tmp & or_18_cse;
  assign and_56_nl = or_tmp_2 & or_620_cse & mux_343_cse;
  assign mux_tmp_11 = MUX_s_1_2_2(and_58_nl, and_56_nl, main_stage_0_2);
  assign nand_83_nl = ~(O_mac_irrel_at_max_sva & mux_tmp_11);
  assign nand_84_nl = ~(if_for_if_for_and_26_tmp & mux_tmp_11);
  assign mux_345_nl = MUX_s_1_2_2(nand_83_nl, nand_84_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign and_dcpl = ~(mux_345_nl | flags_top_1_1_sva);
  assign and_tmp_14 = or_620_cse & or_tmp_10;
  assign and_64_nl = mux_124_itm_1 & and_tmp_14;
  assign and_63_nl = O_wr_data_rsci_ivld_mxwt & and_tmp_14;
  assign mux_346_cse = MUX_s_1_2_2(and_64_nl, and_63_nl, land_9_lpi_1_dfm_1_1);
  assign mux_tmp_14 = MUX_s_1_2_2(mux_346_cse, and_tmp_14, or_1_cse);
  assign nor_tmp_8 = if_for_if_for_and_26_tmp & flags_top_1_1_sva;
  assign not_tmp_8 = ~((if_6_if_3_acc_tmp[0]) & mux_343_cse);
  assign not_tmp_9 = ~(W_irrel_cnt_sva_0 & mux_343_cse);
  assign and_75_nl = mux_124_itm_1 & or_620_cse;
  assign and_74_nl = O_wr_data_rsci_ivld_mxwt & or_620_cse;
  assign mux_356_nl = MUX_s_1_2_2(and_75_nl, and_74_nl, land_9_lpi_1_dfm_1_1);
  assign mux_tmp_24 = MUX_s_1_2_2(mux_356_nl, or_620_cse, or_1_cse);
  assign not_tmp_14 = ~((if_6_if_1_acc_tmp[0]) & mux_tmp_24);
  assign not_tmp_15 = ~(I_irrel_cnt_sva_0 & mux_tmp_24);
  assign and_92_nl = O_mac_irrel_at_max_sva & mux_tmp_14;
  assign and_91_nl = if_for_if_for_and_26_tmp & mux_tmp_14;
  assign mux_tmp_34 = MUX_s_1_2_2(and_92_nl, and_91_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign or_tmp_51 = (~ or_tmp_10) | flags_top_1_1_sva;
  assign nand_14_nl = ~(mux_124_itm_1 & (~ or_tmp_51));
  assign nand_13_nl = ~(O_wr_data_rsci_ivld_mxwt & (~ or_tmp_51));
  assign mux_368_nl = MUX_s_1_2_2(nand_14_nl, nand_13_nl, land_9_lpi_1_dfm_1_1);
  assign mux_369_nl = MUX_s_1_2_2(mux_368_nl, or_tmp_51, or_1_cse);
  assign and_306_cse = or_620_cse & (~ mux_369_nl);
  assign nor_tmp_25 = if_for_if_for_and_26_tmp & oif_2_unequal_tmp;
  assign and_tmp_40 = ((~ or_1_cse) | (~ oif_1_unequal_tmp) | flags_top_1_1_sva)
      & or_18_cse;
  assign nor_tmp_26 = O_mac_irrel_at_max_sva & oif_2_unequal_tmp;
  assign or_dcpl_11 = (~ O_mac_irrel_at_max_sva_dfm_mx0) | flags_top_1_1_sva;
  assign nand_78_cse = ~(or_620_cse & mux_343_cse);
  assign and_305_nl = oif_2_unequal_tmp & (~((~ or_1_cse) | (~ oif_1_unequal_tmp)
      | (skid_buf_top_cnt_sva!=2'b00)));
  assign nor_208_nl = ~((mux1h_7_tmp!=2'b00) | nand_78_cse);
  assign not_tmp_25 = MUX_s_1_2_2(and_305_nl, nor_208_nl, main_stage_0_2);
  assign or_tmp_73 = (~((~ or_1_cse) | (~ oif_1_unequal_tmp) | flags_top_1_1_sva))
      | (skid_buf_top_cnt_sva!=2'b00);
  assign or_dcpl_14 = (mux_188_tmp!=2'b00);
  assign nor_tmp_39 = ~(flags_wr_zero_guard_sva | (~ wr_data_zero_guard_rsci_ivld_mxwt));
  assign nor_tmp_43 = oif_2_unequal_tmp & oif_1_unequal_tmp;
  assign mux_396_cse = MUX_s_1_2_2(nor_tmp_43, and_tmp_14, main_stage_0_2);
  assign or_569_cse = (~ if_6_aif_equal_tmp) | (~ libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_21)
      | (if_6_if_6_mux1h_tmp!=5'b00000);
  assign or_tmp_93 = land_lpi_1_dfm_1 | (~(or_569_cse & main_stage_0_2 & or_620_cse
      & if_6_else_if_equal_tmp & mux_342_cse));
  assign nor_203_nl = ~(and_526_cse | or_tmp_93);
  assign nor_204_nl = ~(nor_tmp_8 | or_tmp_93);
  assign mux_399_nl = MUX_s_1_2_2(nor_203_nl, nor_204_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign or_119_nl = and_526_cse | (~ if_6_aif_equal_tmp) | (~ libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_21)
      | (if_6_if_6_mux1h_tmp!=5'b00000) | (~ mux_396_cse);
  assign or_117_nl = nor_tmp_8 | (~ if_6_aif_equal_tmp) | (~ libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_21)
      | (if_6_if_6_mux1h_tmp!=5'b00000) | (~ mux_396_cse);
  assign mux_397_nl = MUX_s_1_2_2(or_119_nl, or_117_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign mux_tmp_67 = MUX_s_1_2_2(mux_399_nl, mux_397_nl, O_data_vld_sva);
  assign or_tmp_96 = wr_data_zero_guard_rsci_idat_mxwt | mux_tmp_67;
  assign or_tmp_97 = skid_buf_wr_zero_guard_regs_0_sva_dfm_1 | mux_tmp_67;
  assign or_tmp_98 = skid_buf_wr_zero_guard_regs_1_sva_dfm_1 | mux_tmp_67;
  assign mux_404_tmp = MUX_s_1_2_2(or_tmp_97, or_tmp_98, skid_buf_wr_zero_guard_rd_ptr_sva);
  assign mux_402_nl = MUX_s_1_2_2(or_tmp_96, or_tmp_98, skid_buf_wr_zero_guard_rd_ptr_sva);
  assign mux_401_nl = MUX_s_1_2_2(or_tmp_97, or_tmp_96, skid_buf_wr_zero_guard_rd_ptr_sva);
  assign mux_403_nl = MUX_s_1_2_2(mux_402_nl, mux_401_nl, skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_405_cse = MUX_s_1_2_2(mux_404_tmp, mux_403_nl, nor_tmp_39);
  assign and_dcpl_19 = (~ mux_405_cse) & or_dcpl_14 & aif_7_equal_tmp;
  assign or_dcpl_19 = (~ W_wr_data_rsci_ivld_mxwt) | W_data_vld_sva_dfm_1_1;
  assign or_dcpl_21 = or_dcpl_19 | (~ main_stage_0_2) | (W_wr_pntr_sva!=5'b00000);
  assign or_dcpl_22 = (W_wr_pntr_sva[0]) | (W_wr_pntr_sva[2]);
  assign or_dcpl_23 = or_dcpl_22 | (W_wr_pntr_sva[4]);
  assign or_dcpl_25 = or_dcpl_19 | (W_wr_pntr_sva[3]) | (W_wr_pntr_sva[1]);
  assign or_dcpl_27 = (~ (W_wr_pntr_sva[0])) | (W_wr_pntr_sva[2]);
  assign or_dcpl_28 = or_dcpl_27 | (W_wr_pntr_sva[4]);
  assign or_dcpl_29 = or_dcpl_25 | or_dcpl_28;
  assign or_dcpl_31 = or_dcpl_19 | (W_wr_pntr_sva[3]) | (~ (W_wr_pntr_sva[1]));
  assign or_dcpl_32 = or_dcpl_31 | or_dcpl_23;
  assign or_dcpl_33 = or_dcpl_31 | or_dcpl_28;
  assign or_dcpl_34 = (W_wr_pntr_sva[0]) | (~ (W_wr_pntr_sva[2]));
  assign or_dcpl_35 = or_dcpl_34 | (W_wr_pntr_sva[4]);
  assign or_dcpl_36 = or_dcpl_25 | or_dcpl_35;
  assign or_dcpl_37 = ~((W_wr_pntr_sva[0]) & (W_wr_pntr_sva[2]));
  assign or_dcpl_38 = or_dcpl_37 | (W_wr_pntr_sva[4]);
  assign or_dcpl_39 = or_dcpl_25 | or_dcpl_38;
  assign or_dcpl_40 = or_dcpl_31 | or_dcpl_35;
  assign or_dcpl_41 = or_dcpl_31 | or_dcpl_38;
  assign or_dcpl_43 = or_dcpl_19 | (~ (W_wr_pntr_sva[3])) | (W_wr_pntr_sva[1]);
  assign or_dcpl_44 = or_dcpl_43 | or_dcpl_23;
  assign or_dcpl_45 = or_dcpl_43 | or_dcpl_28;
  assign or_dcpl_47 = or_dcpl_19 | (~ (W_wr_pntr_sva[3])) | (~ (W_wr_pntr_sva[1]));
  assign or_dcpl_48 = or_dcpl_47 | or_dcpl_23;
  assign or_dcpl_49 = or_dcpl_47 | or_dcpl_28;
  assign or_dcpl_50 = or_dcpl_43 | or_dcpl_35;
  assign or_dcpl_51 = or_dcpl_43 | or_dcpl_38;
  assign or_dcpl_52 = or_dcpl_47 | or_dcpl_35;
  assign or_dcpl_53 = or_dcpl_47 | or_dcpl_38;
  assign or_dcpl_54 = or_dcpl_22 | (~ (W_wr_pntr_sva[4]));
  assign or_dcpl_55 = or_dcpl_25 | or_dcpl_54;
  assign or_dcpl_56 = or_dcpl_27 | (~ (W_wr_pntr_sva[4]));
  assign or_dcpl_57 = or_dcpl_25 | or_dcpl_56;
  assign or_dcpl_58 = or_dcpl_31 | or_dcpl_54;
  assign or_dcpl_59 = or_dcpl_31 | or_dcpl_56;
  assign or_dcpl_60 = or_dcpl_34 | (~ (W_wr_pntr_sva[4]));
  assign or_dcpl_61 = or_dcpl_25 | or_dcpl_60;
  assign or_dcpl_62 = or_dcpl_37 | (~ (W_wr_pntr_sva[4]));
  assign or_dcpl_63 = or_dcpl_25 | or_dcpl_62;
  assign or_dcpl_64 = or_dcpl_31 | or_dcpl_60;
  assign or_dcpl_65 = or_dcpl_31 | or_dcpl_62;
  assign or_dcpl_66 = or_dcpl_43 | or_dcpl_54;
  assign or_dcpl_67 = or_dcpl_43 | or_dcpl_56;
  assign or_dcpl_68 = or_dcpl_47 | or_dcpl_54;
  assign or_dcpl_69 = or_dcpl_47 | or_dcpl_56;
  assign or_dcpl_70 = or_dcpl_43 | or_dcpl_60;
  assign or_dcpl_71 = or_dcpl_43 | or_dcpl_62;
  assign or_dcpl_72 = or_dcpl_47 | or_dcpl_60;
  assign or_dcpl_73 = or_dcpl_47 | or_dcpl_62;
  assign nand_75_nl = ~(oif_2_unequal_tmp & or_1_cse & oif_1_unequal_tmp);
  assign not_tmp_47 = MUX_s_1_2_2(nand_75_nl, nand_78_cse, main_stage_0_2);
  assign or_192_nl = and_526_cse | not_tmp_47;
  assign or_191_nl = nor_tmp_8 | not_tmp_47;
  assign mux_tmp_76 = MUX_s_1_2_2(or_192_nl, or_191_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign or_dcpl_78 = (~ I_wr_data_rsci_ivld_mxwt) | I_data_vld_sva_dfm_1_1;
  assign or_dcpl_80 = or_dcpl_78 | (~ main_stage_0_2) | (I_wr_pntr_sva!=5'b00000);
  assign or_dcpl_81 = (I_wr_pntr_sva[1]) | (I_wr_pntr_sva[3]);
  assign or_dcpl_82 = or_dcpl_81 | (I_wr_pntr_sva[4]);
  assign or_dcpl_84 = or_dcpl_78 | (I_wr_pntr_sva[0]) | (I_wr_pntr_sva[2]);
  assign or_dcpl_87 = or_dcpl_78 | (~ (I_wr_pntr_sva[0])) | (I_wr_pntr_sva[2]);
  assign or_dcpl_88 = or_dcpl_87 | or_dcpl_82;
  assign or_dcpl_89 = (~ (I_wr_pntr_sva[1])) | (I_wr_pntr_sva[3]);
  assign or_dcpl_90 = or_dcpl_89 | (I_wr_pntr_sva[4]);
  assign or_dcpl_91 = or_dcpl_84 | or_dcpl_90;
  assign or_dcpl_92 = or_dcpl_87 | or_dcpl_90;
  assign or_dcpl_94 = or_dcpl_78 | (I_wr_pntr_sva[0]) | (~ (I_wr_pntr_sva[2]));
  assign or_dcpl_95 = or_dcpl_94 | or_dcpl_82;
  assign or_dcpl_97 = or_dcpl_78 | (~ (I_wr_pntr_sva[0])) | (~ (I_wr_pntr_sva[2]));
  assign or_dcpl_98 = or_dcpl_97 | or_dcpl_82;
  assign or_dcpl_99 = or_dcpl_94 | or_dcpl_90;
  assign or_dcpl_100 = or_dcpl_97 | or_dcpl_90;
  assign or_dcpl_101 = (I_wr_pntr_sva[1]) | (~ (I_wr_pntr_sva[3]));
  assign or_dcpl_102 = or_dcpl_101 | (I_wr_pntr_sva[4]);
  assign or_dcpl_103 = or_dcpl_84 | or_dcpl_102;
  assign or_dcpl_104 = or_dcpl_87 | or_dcpl_102;
  assign or_dcpl_105 = ~((I_wr_pntr_sva[1]) & (I_wr_pntr_sva[3]));
  assign or_dcpl_106 = or_dcpl_105 | (I_wr_pntr_sva[4]);
  assign or_dcpl_107 = or_dcpl_84 | or_dcpl_106;
  assign or_dcpl_108 = or_dcpl_87 | or_dcpl_106;
  assign or_dcpl_109 = or_dcpl_94 | or_dcpl_102;
  assign or_dcpl_110 = or_dcpl_97 | or_dcpl_102;
  assign or_dcpl_111 = or_dcpl_94 | or_dcpl_106;
  assign or_dcpl_112 = or_dcpl_97 | or_dcpl_106;
  assign or_dcpl_113 = or_dcpl_81 | (~ (I_wr_pntr_sva[4]));
  assign or_dcpl_114 = or_dcpl_84 | or_dcpl_113;
  assign or_dcpl_115 = or_dcpl_87 | or_dcpl_113;
  assign or_dcpl_116 = or_dcpl_89 | (~ (I_wr_pntr_sva[4]));
  assign or_dcpl_117 = or_dcpl_84 | or_dcpl_116;
  assign or_dcpl_118 = or_dcpl_87 | or_dcpl_116;
  assign or_dcpl_119 = or_dcpl_94 | or_dcpl_113;
  assign or_dcpl_120 = or_dcpl_97 | or_dcpl_113;
  assign or_dcpl_121 = or_dcpl_94 | or_dcpl_116;
  assign or_dcpl_122 = or_dcpl_97 | or_dcpl_116;
  assign or_dcpl_123 = or_dcpl_101 | (~ (I_wr_pntr_sva[4]));
  assign or_dcpl_124 = or_dcpl_84 | or_dcpl_123;
  assign or_dcpl_125 = or_dcpl_87 | or_dcpl_123;
  assign or_dcpl_126 = or_dcpl_105 | (~ (I_wr_pntr_sva[4]));
  assign or_dcpl_127 = or_dcpl_84 | or_dcpl_126;
  assign or_dcpl_128 = or_dcpl_87 | or_dcpl_126;
  assign or_dcpl_129 = or_dcpl_94 | or_dcpl_123;
  assign or_dcpl_130 = or_dcpl_97 | or_dcpl_123;
  assign or_dcpl_131 = or_dcpl_94 | or_dcpl_126;
  assign or_dcpl_132 = or_dcpl_97 | or_dcpl_126;
  assign and_tmp_56 = flags_top_1_1_sva & O_mac_irrel_at_max_sva_dfm_mx0;
  assign or_tmp_105 = and_541_cse | oif_2_unequal_tmp;
  assign nand_31_nl = ~(or_tmp_105 & (~ and_tmp_56));
  assign mux_tmp_77 = MUX_s_1_2_2(nand_31_nl, and_tmp_56, W_data_vld_sva_dfm_1_1);
  assign or_tmp_106 = and_295_cse | oif_1_unequal_tmp;
  assign nand_32_nl = ~(or_tmp_106 & (~ mux_tmp_77));
  assign mux_tmp_78 = MUX_s_1_2_2(nand_32_nl, mux_tmp_77, I_data_vld_sva_dfm_1_1);
  assign and_tmp_57 = O_data_vld_sva & mux_tmp_78;
  assign nand_34_nl = ~(or_tmp_105 & oif_unequal_tmp & (~ and_tmp_56));
  assign nand_33_nl = ~(oif_unequal_tmp & (~ and_tmp_56));
  assign mux_tmp_79 = MUX_s_1_2_2(nand_34_nl, nand_33_nl, W_data_vld_sva_dfm_1_1);
  assign nand_35_nl = ~(or_tmp_106 & (~ mux_tmp_79));
  assign mux_413_nl = MUX_s_1_2_2(nand_35_nl, mux_tmp_79, I_data_vld_sva_dfm_1_1);
  assign mux_414_nl = MUX_s_1_2_2(mux_413_nl, mux_tmp_78, O_data_vld_sva);
  assign not_tmp_56 = ~(land_lpi_1_dfm_1 | mux_414_nl);
  assign mux_416_nl = MUX_s_1_2_2(not_tmp_56, and_tmp_57, mux_124_itm_1);
  assign mux_415_nl = MUX_s_1_2_2(not_tmp_56, and_tmp_57, O_wr_data_rsci_ivld_mxwt);
  assign mux_tmp_84 = MUX_s_1_2_2(mux_416_nl, mux_415_nl, land_9_lpi_1_dfm_1_1);
  assign or_dcpl_136 = (O_mac_pntr_sva[1:0]!=2'b00);
  assign or_dcpl_137 = (O_mac_pntr_sva[3:2]!=2'b00);
  assign or_dcpl_138 = or_dcpl_137 | or_dcpl_136;
  assign or_dcpl_139 = O_mac_irrel_at_max_sva_dfm_mx0 | (O_mac_pntr_sva[4]);
  assign nor_tmp_65 = if_9_if_equal_1_tmp & I_wr_data_rsci_ivld_mxwt & main_stage_0_2;
  assign mux_tmp_89 = MUX_s_1_2_2(nor_tmp_65, main_stage_0_2, or_tmp_5);
  assign and_128_nl = mux_124_itm_1 & mux_tmp_89;
  assign and_127_nl = O_wr_data_rsci_ivld_mxwt & mux_tmp_89;
  assign mux_tmp_91 = MUX_s_1_2_2(and_128_nl, and_127_nl, land_9_lpi_1_dfm_1_1);
  assign and_129_nl = or_558_cse & mux_tmp_91;
  assign mux_425_nl = MUX_s_1_2_2(and_129_nl, mux_tmp_91, oif_2_unequal_tmp);
  assign and_126_nl = or_558_cse & mux_tmp_89;
  assign mux_421_nl = MUX_s_1_2_2(nor_tmp_65, main_stage_0_2, I_data_vld_sva_dfm_1_1);
  assign or_267_nl = oif_1_unequal_tmp | mux_421_nl;
  assign mux_423_nl = MUX_s_1_2_2(and_126_nl, or_267_nl, oif_2_unequal_tmp);
  assign mux_426_itm = MUX_s_1_2_2(mux_425_nl, mux_423_nl, or_1_cse);
  assign or_dcpl_142 = (O_mac_pntr_sva[1:0]!=2'b01);
  assign or_dcpl_143 = or_dcpl_137 | or_dcpl_142;
  assign or_dcpl_146 = (O_mac_pntr_sva[1:0]!=2'b10);
  assign or_dcpl_147 = or_dcpl_137 | or_dcpl_146;
  assign or_dcpl_150 = ~((O_mac_pntr_sva[1:0]==2'b11));
  assign or_dcpl_151 = or_dcpl_137 | or_dcpl_150;
  assign or_dcpl_154 = (O_mac_pntr_sva[3:2]!=2'b01);
  assign or_dcpl_155 = or_dcpl_154 | or_dcpl_136;
  assign or_dcpl_158 = or_dcpl_154 | or_dcpl_142;
  assign or_dcpl_161 = or_dcpl_154 | or_dcpl_146;
  assign or_dcpl_164 = or_dcpl_154 | or_dcpl_150;
  assign or_dcpl_167 = (O_mac_pntr_sva[3:2]!=2'b10);
  assign or_dcpl_168 = or_dcpl_167 | or_dcpl_136;
  assign or_dcpl_171 = or_dcpl_167 | or_dcpl_142;
  assign or_dcpl_174 = or_dcpl_167 | or_dcpl_146;
  assign or_dcpl_177 = or_dcpl_167 | or_dcpl_150;
  assign or_dcpl_180 = ~((O_mac_pntr_sva[3:2]==2'b11));
  assign or_dcpl_181 = or_dcpl_180 | or_dcpl_136;
  assign or_dcpl_184 = or_dcpl_180 | or_dcpl_142;
  assign or_dcpl_187 = or_dcpl_180 | or_dcpl_146;
  assign or_dcpl_190 = or_dcpl_180 | or_dcpl_150;
  assign or_dcpl_193 = O_mac_irrel_at_max_sva_dfm_mx0 | (~ (O_mac_pntr_sva[4]));
  assign or_dcpl_226 = ~(main_stage_0_2 & or_svs_1);
  assign nor_201_nl = ~(skid_buf_top_wr_ptr_sva_1 | skid_buf_top_wr_ptr_sva_0);
  assign mux_tmp_94 = MUX_s_1_2_2(nor_201_nl, skid_buf_top_push_nor_psp, if_5_and_svs_1);
  assign nor_200_nl = ~(skid_buf_top_wr_ptr_sva_1 | (~ skid_buf_top_wr_ptr_sva_0));
  assign mux_tmp_96 = MUX_s_1_2_2(nor_200_nl, skid_buf_top_push_and_psp, if_5_and_svs_1);
  assign nor_199_nl = ~((~ skid_buf_top_wr_ptr_sva_1) | skid_buf_top_wr_ptr_sva_0);
  assign mux_tmp_98 = MUX_s_1_2_2(nor_199_nl, skid_buf_top_push_and_1_psp, if_5_and_svs_1);
  assign or_dcpl_237 = ~(or_dcpl_14 & aif_7_equal_tmp);
  assign or_tmp_143 = land_lpi_1_dfm_1 | (~(or_569_cse & if_6_else_if_equal_tmp &
      mux_346_cse));
  assign nor_195_nl = ~(and_526_cse | or_tmp_143);
  assign nor_196_nl = ~(nor_tmp_8 | or_tmp_143);
  assign mux_445_nl = MUX_s_1_2_2(nor_195_nl, nor_196_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign or_394_nl = and_526_cse | (~ if_6_aif_equal_tmp) | (~ libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_21)
      | (if_6_if_6_mux1h_tmp!=5'b00000) | (~ and_tmp_14);
  assign or_392_nl = nor_tmp_8 | (~ if_6_aif_equal_tmp) | (~ libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_21)
      | (if_6_if_6_mux1h_tmp!=5'b00000) | (~ and_tmp_14);
  assign mux_443_nl = MUX_s_1_2_2(or_394_nl, or_392_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign mux_tmp_113 = MUX_s_1_2_2(mux_445_nl, mux_443_nl, O_data_vld_sva);
  assign or_399_cse = wr_data_zero_guard_rsci_idat_mxwt | mux_tmp_113;
  assign or_400_cse = skid_buf_wr_zero_guard_regs_0_sva_dfm_1 | mux_tmp_113;
  assign or_401_cse = skid_buf_wr_zero_guard_regs_1_sva_dfm_1 | mux_tmp_113;
  assign or_tmp_162 = (~ wr_data_zero_guard_rsci_ivld_mxwt) | flags_wr_zero_guard_sva;
  assign not_tmp_93 = ~(or_620_cse & or_tmp_10);
  assign or_422_nl = O_mac_irrel_at_max_sva | not_tmp_93;
  assign or_421_nl = if_for_if_for_and_26_tmp | not_tmp_93;
  assign mux_461_nl = MUX_s_1_2_2(or_422_nl, or_421_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign mux_tmp_129 = MUX_s_1_2_2(not_tmp_93, mux_461_nl, flags_top_1_1_sva);
  assign nor_110_cse = ~((~ libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_21)
      | (if_6_if_6_mux1h_tmp!=5'b00000) | (~ if_6_aif_equal_tmp));
  assign nor_191_nl = ~(O_mac_irrel_at_max_sva | (~ nor_tmp_43));
  assign nor_192_nl = ~(if_for_if_for_and_26_tmp | (~ nor_tmp_43));
  assign mux_463_nl = MUX_s_1_2_2(nor_191_nl, nor_192_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign mux_464_nl = MUX_s_1_2_2(nor_tmp_43, mux_463_nl, flags_top_1_1_sva);
  assign mux_465_nl = MUX_s_1_2_2(mux_464_nl, (~ mux_tmp_129), main_stage_0_2);
  assign nand_tmp_25 = ~(nor_110_cse & mux_465_nl);
  assign and_299_nl = or_569_cse & main_stage_0_2 & (~ mux_tmp_129);
  assign mux_466_nl = MUX_s_1_2_2(and_299_nl, nand_tmp_25, O_data_vld_sva);
  assign nand_tmp_27 = ~(or_dcpl_14 & aif_7_equal_tmp & (~ mux_466_nl));
  assign mux_tmp_134 = MUX_s_1_2_2((~ nand_tmp_27), nand_tmp_27, skid_buf_wr_zero_guard_rd_ptr_sva);
  assign or_tmp_171 = (~ skid_buf_wr_zero_guard_regs_0_sva_dfm_1) | skid_buf_wr_zero_guard_rd_ptr_sva;
  assign nand_tmp_28 = ~(or_tmp_171 & (~ nand_tmp_27));
  assign nor_tmp_110 = skid_buf_wr_zero_guard_regs_1_sva_dfm_1 & skid_buf_wr_zero_guard_rd_ptr_sva;
  assign or_428_nl = nor_tmp_110 | nand_tmp_27;
  assign mux_474_nl = MUX_s_1_2_2(or_428_nl, nand_tmp_28, skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_473_nl = MUX_s_1_2_2(mux_tmp_134, (~ mux_tmp_134), skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_475_nl = MUX_s_1_2_2(mux_474_nl, mux_473_nl, wr_data_zero_guard_rsci_idat_mxwt);
  assign mux_471_nl = MUX_s_1_2_2(nand_tmp_28, (~ mux_tmp_134), skid_buf_wr_zero_guard_regs_1_sva_dfm_1);
  assign mux_469_nl = MUX_s_1_2_2((~ nand_tmp_27), nand_tmp_27, or_tmp_171);
  assign or_425_nl = skid_buf_wr_zero_guard_rd_ptr_sva | nand_tmp_27;
  assign mux_468_nl = MUX_s_1_2_2(or_425_nl, mux_tmp_134, skid_buf_wr_zero_guard_regs_0_sva_dfm_1);
  assign mux_470_nl = MUX_s_1_2_2(mux_469_nl, mux_468_nl, skid_buf_wr_zero_guard_regs_1_sva_dfm_1);
  assign mux_472_nl = MUX_s_1_2_2(mux_471_nl, mux_470_nl, skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_tmp_143 = MUX_s_1_2_2(mux_475_nl, mux_472_nl, or_tmp_162);
  assign nand_tmp_29 = ~(or_dcpl_14 & aif_7_equal_tmp & (~(O_data_vld_sva & nand_tmp_25)));
  assign mux_tmp_144 = MUX_s_1_2_2((~ nand_tmp_29), nand_tmp_29, skid_buf_wr_zero_guard_rd_ptr_sva);
  assign nand_tmp_30 = ~(or_tmp_171 & (~ nand_tmp_29));
  assign or_434_nl = nor_tmp_110 | nand_tmp_29;
  assign mux_484_nl = MUX_s_1_2_2(or_434_nl, nand_tmp_30, skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_483_nl = MUX_s_1_2_2(mux_tmp_144, (~ mux_tmp_144), skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_485_nl = MUX_s_1_2_2(mux_484_nl, mux_483_nl, wr_data_zero_guard_rsci_idat_mxwt);
  assign mux_481_nl = MUX_s_1_2_2(nand_tmp_30, (~ mux_tmp_144), skid_buf_wr_zero_guard_regs_1_sva_dfm_1);
  assign mux_479_nl = MUX_s_1_2_2((~ nand_tmp_29), nand_tmp_29, or_tmp_171);
  assign or_431_nl = skid_buf_wr_zero_guard_rd_ptr_sva | nand_tmp_29;
  assign mux_478_nl = MUX_s_1_2_2(or_431_nl, mux_tmp_144, skid_buf_wr_zero_guard_regs_0_sva_dfm_1);
  assign mux_480_nl = MUX_s_1_2_2(mux_479_nl, mux_478_nl, skid_buf_wr_zero_guard_regs_1_sva_dfm_1);
  assign mux_482_nl = MUX_s_1_2_2(mux_481_nl, mux_480_nl, skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_tmp_153 = MUX_s_1_2_2(mux_485_nl, mux_482_nl, or_tmp_162);
  assign nand_tmp_31 = (~ libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_21)
      | (if_6_if_6_mux1h_tmp!=5'b00000) | (~ if_6_aif_equal_tmp) | mux_tmp_129;
  assign nor_190_nl = ~(nor_110_cse | mux_tmp_129);
  assign mux_493_nl = MUX_s_1_2_2(nor_190_nl, nand_tmp_31, O_data_vld_sva);
  assign nand_tmp_32 = ~(or_dcpl_14 & aif_7_equal_tmp & (~ mux_493_nl));
  assign mux_tmp_161 = MUX_s_1_2_2((~ nand_tmp_32), nand_tmp_32, skid_buf_wr_zero_guard_rd_ptr_sva);
  assign nand_tmp_33 = ~(or_tmp_171 & (~ nand_tmp_32));
  assign or_445_nl = nor_tmp_110 | nand_tmp_32;
  assign mux_501_nl = MUX_s_1_2_2(or_445_nl, nand_tmp_33, skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_500_nl = MUX_s_1_2_2(mux_tmp_161, (~ mux_tmp_161), skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_502_nl = MUX_s_1_2_2(mux_501_nl, mux_500_nl, wr_data_zero_guard_rsci_idat_mxwt);
  assign mux_498_nl = MUX_s_1_2_2(nand_tmp_33, (~ mux_tmp_161), skid_buf_wr_zero_guard_regs_1_sva_dfm_1);
  assign mux_496_nl = MUX_s_1_2_2((~ nand_tmp_32), nand_tmp_32, or_tmp_171);
  assign or_442_nl = skid_buf_wr_zero_guard_rd_ptr_sva | nand_tmp_32;
  assign mux_495_nl = MUX_s_1_2_2(or_442_nl, mux_tmp_161, skid_buf_wr_zero_guard_regs_0_sva_dfm_1);
  assign mux_497_nl = MUX_s_1_2_2(mux_496_nl, mux_495_nl, skid_buf_wr_zero_guard_regs_1_sva_dfm_1);
  assign mux_499_nl = MUX_s_1_2_2(mux_498_nl, mux_497_nl, skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_tmp_170 = MUX_s_1_2_2(mux_502_nl, mux_499_nl, or_tmp_162);
  assign nand_tmp_34 = ~(or_dcpl_14 & aif_7_equal_tmp & (~(O_data_vld_sva & nand_tmp_31)));
  assign mux_tmp_171 = MUX_s_1_2_2((~ nand_tmp_34), nand_tmp_34, skid_buf_wr_zero_guard_rd_ptr_sva);
  assign nand_tmp_35 = ~(or_tmp_171 & (~ nand_tmp_34));
  assign or_451_nl = nor_tmp_110 | nand_tmp_34;
  assign mux_511_nl = MUX_s_1_2_2(or_451_nl, nand_tmp_35, skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_510_nl = MUX_s_1_2_2(mux_tmp_171, (~ mux_tmp_171), skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_512_nl = MUX_s_1_2_2(mux_511_nl, mux_510_nl, wr_data_zero_guard_rsci_idat_mxwt);
  assign mux_508_nl = MUX_s_1_2_2(nand_tmp_35, (~ mux_tmp_171), skid_buf_wr_zero_guard_regs_1_sva_dfm_1);
  assign mux_506_nl = MUX_s_1_2_2((~ nand_tmp_34), nand_tmp_34, or_tmp_171);
  assign or_448_nl = skid_buf_wr_zero_guard_rd_ptr_sva | nand_tmp_34;
  assign mux_505_nl = MUX_s_1_2_2(or_448_nl, mux_tmp_171, skid_buf_wr_zero_guard_regs_0_sva_dfm_1);
  assign mux_507_nl = MUX_s_1_2_2(mux_506_nl, mux_505_nl, skid_buf_wr_zero_guard_regs_1_sva_dfm_1);
  assign mux_509_nl = MUX_s_1_2_2(mux_508_nl, mux_507_nl, skid_buf_wr_zero_guard_wr_ptr_sva);
  assign mux_tmp_180 = MUX_s_1_2_2(mux_512_nl, mux_509_nl, or_tmp_162);
  assign or_tmp_200 = or_620_cse | or_557_cse;
  assign mux_520_nl = MUX_s_1_2_2(or_557_cse, or_tmp_200, mux_124_itm_1);
  assign mux_519_nl = MUX_s_1_2_2(or_557_cse, or_tmp_200, O_wr_data_rsci_ivld_mxwt);
  assign mux_521_nl = MUX_s_1_2_2(mux_520_nl, mux_519_nl, land_9_lpi_1_dfm_1_1);
  assign and_153_nl = main_stage_0_2 & mux_521_nl;
  assign mux_518_nl = MUX_s_1_2_2(oif_2_unequal_tmp, or_tmp_200, main_stage_0_2);
  assign mux_tmp_189 = MUX_s_1_2_2(and_153_nl, mux_518_nl, or_1_cse);
  assign and_tmp_80 = main_stage_0_2 & or_557_cse;
  assign or_tmp_204 = or_tmp_10 | or_558_cse;
  assign mux_532_nl = MUX_s_1_2_2(or_558_cse, or_tmp_204, mux_124_itm_1);
  assign mux_531_nl = MUX_s_1_2_2(or_558_cse, or_tmp_204, O_wr_data_rsci_ivld_mxwt);
  assign mux_533_nl = MUX_s_1_2_2(mux_532_nl, mux_531_nl, land_9_lpi_1_dfm_1_1);
  assign mux_534_nl = MUX_s_1_2_2(mux_533_nl, or_tmp_204, or_1_cse);
  assign mux_tmp_202 = MUX_s_1_2_2(and_544_cse, mux_534_nl, main_stage_0_2);
  assign and_tmp_81 = main_stage_0_2 & or_558_cse;
  assign or_dcpl_246 = (~ skid_buf_wr_zero_guard_wr_ptr_sva) | flags_wr_zero_guard_sva
      | (~ wr_data_zero_guard_rsci_ivld_mxwt);
  assign or_dcpl_248 = skid_buf_wr_zero_guard_wr_ptr_sva | flags_wr_zero_guard_sva
      | (~ wr_data_zero_guard_rsci_ivld_mxwt);
  assign and_tmp_93 = nor_tmp_65 & or_tmp_2;
  assign mux_tmp_224 = MUX_s_1_2_2(and_tmp_93, and_tmp, or_tmp_5);
  assign and_171_nl = mux_124_itm_1 & mux_tmp_224;
  assign and_170_nl = O_wr_data_rsci_ivld_mxwt & mux_tmp_224;
  assign mux_tmp_226 = MUX_s_1_2_2(and_171_nl, and_170_nl, land_9_lpi_1_dfm_1_1);
  assign and_296_nl = mux_124_itm_1 & main_stage_0_2;
  assign and_297_nl = O_wr_data_rsci_ivld_mxwt & main_stage_0_2;
  assign mux_tmp_231 = MUX_s_1_2_2(and_296_nl, and_297_nl, land_9_lpi_1_dfm_1_1);
  assign mux_tmp_232 = MUX_s_1_2_2(mux_tmp_231, main_stage_0_2, oif_unequal_tmp);
  assign and_tmp_98 = and_295_cse & mux_tmp_232;
  assign and_175_nl = W_data_vld_sva_dfm_1_1 & if_9_if_equal_1_tmp & I_wr_data_rsci_ivld_mxwt
      & mux_tmp_232;
  assign and_174_nl = W_data_vld_sva_dfm_1_1 & mux_tmp_232;
  assign mux_569_nl = MUX_s_1_2_2(and_175_nl, and_174_nl, or_tmp_5);
  assign mux_568_nl = MUX_s_1_2_2(and_tmp_98, mux_tmp_232, or_tmp_5);
  assign mux_570_nl = MUX_s_1_2_2(mux_569_nl, mux_568_nl, and_541_cse);
  assign mux_566_nl = MUX_s_1_2_2(and_tmp_98, mux_tmp_232, I_data_vld_sva_dfm_1_1);
  assign or_493_nl = oif_unequal_tmp | mux_tmp_231;
  assign mux_567_nl = MUX_s_1_2_2(mux_566_nl, or_493_nl, oif_1_unequal_tmp);
  assign mux_571_itm = MUX_s_1_2_2(mux_570_nl, mux_567_nl, oif_2_unequal_tmp);
  assign nor_188_nl = ~(and_526_cse | (~ mux_571_itm));
  assign nor_189_nl = ~(nor_tmp_8 | (~ mux_571_itm));
  assign mux_572_nl = MUX_s_1_2_2(nor_188_nl, nor_189_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign and_dcpl_28 = ~(mux_572_nl | O_data_vld_sva);
  assign or_tmp_242 = and_dcpl_19 & (fsm_output[1]);
  assign O_rd_data_rsci_idat_mx0c0 = (and_dcpl & (fsm_output[1])) | (mux_tmp_34 &
      or_tmp_2 & (~ flags_top_1_1_sva) & main_stage_0_2);
  assign mux_372_nl = MUX_s_1_2_2(or_18_cse, and_tmp_40, nor_tmp_26);
  assign mux_371_nl = MUX_s_1_2_2(or_18_cse, and_tmp_40, nor_tmp_25);
  assign mux_373_nl = MUX_s_1_2_2(mux_372_nl, mux_371_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign nand_17_nl = ~(O_mac_irrel_at_max_sva & and_306_cse);
  assign nand_16_nl = ~(if_for_if_for_and_26_tmp & and_306_cse);
  assign mux_370_nl = MUX_s_1_2_2(nand_17_nl, nand_16_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign and_95_nl = or_tmp_2 & mux_370_nl;
  assign mux_374_nl = MUX_s_1_2_2(mux_373_nl, and_95_nl, main_stage_0_2);
  assign O_rd_data_rsci_idat_mx0c1 = (mux_374_nl & (fsm_output[1])) | (((~ mux_tmp_14)
      | or_dcpl_11) & or_tmp_2 & main_stage_0_2);
  assign nand_57_nl = ~(O_mac_irrel_at_max_sva & not_tmp_25);
  assign nand_58_nl = ~(if_for_if_for_and_26_tmp & not_tmp_25);
  assign mux_381_nl = MUX_s_1_2_2(nand_57_nl, nand_58_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign O_rd_data_rsci_idat_mx0c2 = ((~(mux_381_nl | flags_top_1_1_sva)) & (fsm_output[1]))
      | (mux_tmp_34 & (~ flags_top_1_1_sva) & (mux1h_7_tmp==2'b00) & main_stage_0_2);
  assign O_data_vld_sva_mx0c1 = ((mux_405_cse | or_dcpl_237) & (fsm_output[1])) |
      ((mux_460_cse | or_dcpl_237) & main_stage_0_2);
  assign nor_138_nl = ~(and_526_cse | (I_irrel_cnt_sva_4_1!=4'b0000) | (~ I_irrel_cnt_sva_0));
  assign mux_527_nl = MUX_s_1_2_2(and_tmp_80, mux_tmp_189, nor_138_nl);
  assign nor_136_nl = ~(and_526_cse | (if_6_if_1_acc_tmp!=5'b00001));
  assign mux_526_nl = MUX_s_1_2_2(and_tmp_80, mux_tmp_189, nor_136_nl);
  assign mux_528_nl = MUX_s_1_2_2(mux_527_nl, mux_526_nl, I_mac_irrel_at_maxBuf_sva);
  assign nor_134_nl = ~(nor_tmp_8 | (I_irrel_cnt_sva_4_1!=4'b0000) | (~ I_irrel_cnt_sva_0));
  assign mux_524_nl = MUX_s_1_2_2(and_tmp_80, mux_tmp_189, nor_134_nl);
  assign nor_130_nl = ~(nor_tmp_8 | (if_6_if_1_acc_tmp!=5'b00001));
  assign mux_523_nl = MUX_s_1_2_2(and_tmp_80, mux_tmp_189, nor_130_nl);
  assign mux_525_nl = MUX_s_1_2_2(mux_524_nl, mux_523_nl, if_for_if_for_and_27_tmp);
  assign mux_529_nl = MUX_s_1_2_2(mux_528_nl, mux_525_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign mux_530_itm = MUX_s_1_2_2(and_tmp_80, mux_529_nl, oif_1_unequal_tmp);
  assign nor_149_nl = ~(and_526_cse | (W_irrel_cnt_sva_4_1!=4'b0000) | (~ W_irrel_cnt_sva_0));
  assign mux_540_nl = MUX_s_1_2_2(and_tmp_81, mux_tmp_202, nor_149_nl);
  assign nor_147_nl = ~(and_526_cse | (if_6_if_3_acc_tmp!=5'b00001));
  assign mux_539_nl = MUX_s_1_2_2(and_tmp_81, mux_tmp_202, nor_147_nl);
  assign mux_541_nl = MUX_s_1_2_2(mux_540_nl, mux_539_nl, W_mac_irrel_at_maxBuf_sva);
  assign nor_145_nl = ~(nor_tmp_8 | (W_irrel_cnt_sva_4_1!=4'b0000) | (~ W_irrel_cnt_sva_0));
  assign mux_537_nl = MUX_s_1_2_2(and_tmp_81, mux_tmp_202, nor_145_nl);
  assign nor_140_nl = ~(nor_tmp_8 | (if_6_if_3_acc_tmp!=5'b00001));
  assign mux_536_nl = MUX_s_1_2_2(and_tmp_81, mux_tmp_202, nor_140_nl);
  assign mux_538_nl = MUX_s_1_2_2(mux_537_nl, mux_536_nl, if_for_if_for_and_28_tmp);
  assign mux_542_nl = MUX_s_1_2_2(mux_541_nl, mux_538_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign mux_543_itm = MUX_s_1_2_2(and_tmp_81, mux_542_nl, oif_2_unequal_tmp);
  assign flags_top_1_1_sva_mx0c1 = (~ main_stage_0_2) & (fsm_output[1]);
  assign or_360_tmp = (~ mux_tmp_94) | or_dcpl_226;
  assign skid_buf_top_peek_and_m1c = (~ skid_buf_top_push_nor_psp_mx0w0) & skid_buf_top_peek_nor_m1c_1;
  assign or_364_tmp = (~ mux_tmp_96) | or_dcpl_226;
  assign skid_buf_top_peek_and_4_m1c = (~ skid_buf_top_push_and_psp_1) & skid_buf_top_peek_and_m1c_2;
  assign or_368_tmp = (~ mux_tmp_98) | or_dcpl_226;
  assign skid_buf_top_peek_and_5_m1c = (~ skid_buf_top_push_and_1_psp_mx0w0) & skid_buf_top_peek_and_m1c_3;
  assign if_5_if_and_3_m1c = skid_buf_top_peek_nor_m1c_1 & O_rd_data_rsci_idat_mx0c1;
  assign if_5_if_and_4_m1c = skid_buf_top_rd_ptr_sva_0_mx1 & (~ skid_buf_top_rd_ptr_sva_1_mx1)
      & O_rd_data_rsci_idat_mx0c1;
  assign if_5_if_and_5_m1c = skid_buf_top_rd_ptr_sva_1_mx1 & (~ skid_buf_top_rd_ptr_sva_0_mx1)
      & O_rd_data_rsci_idat_mx0c1;
  assign and_331_cse = nand_73_cse & (fsm_output[1]);
  assign and_dcpl_34 = or_svs_1 & main_stage_0_2;
  assign or_dcpl = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1_1
      | if_5_and_svs_1;
  assign mux_585_nl = MUX_s_1_2_2((~ O_rd_data_rsci_irdy_mxwt), O_rd_data_rsci_irdy_mxwt,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1_1);
  assign or_tmp_299 = if_5_and_svs_1 | mux_585_nl;
  assign or_tmp_300 = oif_2_unequal_tmp | W_data_vld_sva_dfm_1_1;
  assign or_756_cse = (O_instr_in_rsci_idat_mxwt[24:0]!=25'b0000100001000010000100001);
  assign not_tmp_156 = ~(or_756_cse & reg_W_instr_in_rsci_oswt_cse_1);
  assign or_598_cse = (z_out_3!=2'b00);
  assign nand_tmp = ~(or_598_cse & not_tmp_156);
  assign or_601_cse = (skid_buf_top_push_1_acc_1_tmp!=2'b00);
  assign or_600_cse = (skid_buf_top_cnt_sva_1_1!=2'b00);
  assign nor_307_nl = ~(O_rd_data_rsci_irdy_mxwt | (or_601_cse & not_tmp_156));
  assign and_365_nl = O_rd_data_rsci_irdy_mxwt & nand_tmp;
  assign mux_587_nl = MUX_s_1_2_2(nor_307_nl, and_365_nl, operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1_1);
  assign nand_96_nl = ~(or_600_cse & not_tmp_156);
  assign mux_586_nl = MUX_s_1_2_2(nand_96_nl, nand_tmp, O_rd_data_rsci_irdy_mxwt);
  assign mux_tmp_245 = MUX_s_1_2_2(mux_587_nl, mux_586_nl, if_5_and_svs_1);
  assign mux_589_nl = MUX_s_1_2_2(or_tmp_299, mux_tmp_245, and_295_cse);
  assign mux_tmp_247 = MUX_s_1_2_2(mux_589_nl, mux_tmp_245, or_tmp_5);
  assign mux_592_nl = MUX_s_1_2_2(or_tmp_299, mux_tmp_247, mux_124_itm_1);
  assign mux_591_nl = MUX_s_1_2_2(or_tmp_299, mux_tmp_247, O_wr_data_rsci_ivld_mxwt);
  assign mux_593_nl = MUX_s_1_2_2(mux_592_nl, mux_591_nl, land_9_lpi_1_dfm_1_1);
  assign mux_tmp_251 = MUX_s_1_2_2(mux_593_nl, mux_tmp_247, or_1_cse);
  assign nor_215_cse = ~((O_instr_in_rsci_idat_mxwt[24:0]!=25'b0000100001000010000100001)
      | (~ O_mac_irrel_at_max_sva) | (~ flags_top_1_1_sva));
  assign and_539_nl = W_mac_irrel_at_maxBuf_sva & nand_129_cse;
  assign nor_304_nl = ~(nor_215_cse | (W_instr_in_rsci_idat_mxwt[24:0]!=25'b0000100001000010000100001));
  assign not_tmp_165 = MUX_s_1_2_2(and_539_nl, nor_304_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign nand_tmp_39 = ~(or_tmp_10 & not_tmp_165);
  assign and_535_nl = I_mac_irrel_at_maxBuf_sva & nand_129_cse;
  assign nor_301_nl = ~(nor_215_cse | (I_instr_in_rsci_idat_mxwt[24:0]!=25'b0000100001000010000100001));
  assign not_tmp_172 = MUX_s_1_2_2(and_535_nl, nor_301_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign nand_tmp_46 = ~(or_tmp_10 & not_tmp_172);
  assign and_dcpl_58 = reg_W_instr_in_rsci_oswt_cse_1 & run_wen;
  assign nor_tmp_182 = or_756_cse & reg_W_instr_in_rsci_oswt_cse_1;
  assign and_tmp_102 = or_tmp_10 & nor_tmp_182;
  assign and_tmp_103 = or_1_cse & aif_equal_tmp & data_zg_sva & nor_tmp_182;
  assign and_tmp_104 = or_tmp_10 & and_tmp_103;
  assign nor_tmp_189 = or_1_cse & aif_equal_tmp & data_zg_sva;
  assign and_tmp_107 = or_tmp_10 & nor_tmp_189;
  assign mux_636_nl = MUX_s_1_2_2(or_601_cse, or_18_cse, operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1_1);
  assign mux_637_nl = MUX_s_1_2_2(mux_636_nl, or_600_cse, if_5_and_svs_1);
  assign mux_635_nl = MUX_s_1_2_2(or_18_cse, or_598_cse, or_dcpl);
  assign mux_638_nl = MUX_s_1_2_2(mux_637_nl, mux_635_nl, O_rd_data_rsci_irdy_mxwt);
  assign mux_tmp_296 = MUX_s_1_2_2(or_18_cse, mux_638_nl, or_svs_1);
  assign not_tmp_191 = nand_129_cse & mux_tmp_296;
  assign not_tmp_193 = ~(nor_tmp_182 | (~ O_mac_irrel_at_max_sva) | flags_top_1_1_sva
      | (~ mux_tmp_296));
  assign and_516_nl = libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_21
      & not_tmp_191;
  assign mux_640_nl = MUX_s_1_2_2(not_tmp_191, mux_tmp_296, reg_W_instr_in_rsci_oswt_cse_1);
  assign and_425_nl = libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_21
      & mux_640_nl;
  assign mux_641_nl = MUX_s_1_2_2(and_516_nl, and_425_nl, or_756_cse);
  assign mux_642_itm = MUX_s_1_2_2(not_tmp_193, mux_641_nl, or_tmp_10);
  assign nor_tmp_217 = (fsm_output[1]) & reg_W_instr_in_rsci_oswt_cse_1;
  assign mux_662_nl = MUX_s_1_2_2((fsm_output[1]), reg_W_instr_in_rsci_oswt_cse_1,
      and_526_cse);
  assign mux_661_nl = MUX_s_1_2_2((fsm_output[1]), nor_tmp_217, and_526_cse);
  assign mux_663_itm = MUX_s_1_2_2(mux_662_nl, mux_661_nl, or_756_cse);
  always @(posedge clk) begin
    if ( rst ) begin
      reg_W_instr_in_rsci_oswt_cse_1 <= 1'b0;
      reg_wr_data_zero_guard_rsci_oswt_cse <= 1'b0;
      reg_W_wr_data_rsci_irdy_run_psct_cse <= 1'b0;
      reg_I_wr_data_rsci_irdy_run_psct_cse <= 1'b0;
      reg_O_rd_data_rsci_ivld_run_psct_cse <= 1'b0;
      reg_O_wr_data_rsci_irdy_run_psct_cse <= 1'b0;
      W_data_vld_sva_dfm_1_1 <= 1'b0;
      I_data_vld_sva_dfm_1_1 <= 1'b0;
      land_9_lpi_1_dfm_1_1 <= 1'b0;
      mac_data_data_sva_dfm_2_1 <= 16'b0000000000000000;
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1_1 <=
          1'b0;
      if_5_and_svs_1 <= 1'b0;
      or_svs_1 <= 1'b0;
      mux_124_itm_1 <= 1'b0;
      data_zg_sva <= 1'b0;
      main_stage_0_2 <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_W_instr_in_rsci_oswt_cse_1 <= ~ (fsm_output[1]);
      reg_wr_data_zero_guard_rsci_oswt_cse <= ~(operator_2_false_5_operator_2_false_5_operator_2_false_5_or_cse
          & (fsm_output[1]));
      reg_W_wr_data_rsci_irdy_run_psct_cse <= (mux_355_nl | (~(or_558_cse & main_stage_0_2)))
          & (fsm_output[1]);
      reg_I_wr_data_rsci_irdy_run_psct_cse <= (mux_360_nl | (~(or_557_cse & main_stage_0_2)))
          & (fsm_output[1]);
      reg_O_rd_data_rsci_ivld_run_psct_cse <= mux_388_nl & (fsm_output[1]);
      reg_O_wr_data_rsci_irdy_run_psct_cse <= or_tmp_242;
      W_data_vld_sva_dfm_1_1 <= MUX_s_1_2_2(if_6_if_6_and_3_nl, W_data_vld_sva_mx0,
          mux_tmp_76);
      I_data_vld_sva_dfm_1_1 <= MUX_s_1_2_2(if_6_if_6_and_nl, I_data_vld_sva_mx0,
          mux_tmp_76);
      land_9_lpi_1_dfm_1_1 <= land_9_lpi_1_dfm_1;
      mac_data_data_sva_dfm_2_1 <= mac_data_data_sva_dfm_3;
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1_1 <=
          operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1;
      if_5_and_svs_1 <= land_5_lpi_1_dfm_1 & operator_2_false_1_operator_2_false_1_operator_2_false_1_or_cse_sva_1;
      or_svs_1 <= land_5_lpi_1_dfm_1 | (skid_buf_top_cnt_sva_mx1!=2'b00);
      mux_124_itm_1 <= MUX_s_1_2_2(if_6_if_6_and_9_nl, O_write_flag_sva_mx0, mux_tmp_76);
      data_zg_sva <= ~((~(mux_123_nl | else_8_land_lpi_1_dfm_mx1)) | land_9_lpi_1_dfm_1);
      main_stage_0_2 <= fsm_output[1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_rd_data_rsci_idat <= 16'b0000000000000000;
    end
    else if ( run_wen & (O_rd_data_rsci_idat_mx0c0 | O_rd_data_rsci_idat_mx0c1 |
        O_rd_data_rsci_idat_mx0c2) ) begin
      O_rd_data_rsci_idat <= MUX1HOT_v_16_5_2(mac_data_data_sva_dfm_2_1, skid_buf_top_regs_data_0_0_sva,
          mac_data_data_sva_dfm_3, skid_buf_top_regs_data_1_0_sva, skid_buf_top_regs_data_2_0_sva,
          {if_5_if_or_nl , if_5_if_or_2_nl , if_5_if_or_3_nl , if_5_if_or_4_nl ,
          if_5_if_or_5_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      flags_wr_zero_guard_sva <= 1'b0;
    end
    else if ( flags_wr_zero_guard_and_cse ) begin
      flags_wr_zero_guard_sva <= operator_2_false_5_operator_2_false_5_operator_2_false_5_or_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_0_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_21) ) begin
      W_mem_0_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_1_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_29) ) begin
      W_mem_1_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_2_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_32) ) begin
      W_mem_2_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_3_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_33) ) begin
      W_mem_3_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_4_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_36) ) begin
      W_mem_4_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_5_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_39) ) begin
      W_mem_5_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_6_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_40) ) begin
      W_mem_6_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_7_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_41) ) begin
      W_mem_7_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_8_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_44) ) begin
      W_mem_8_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_9_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_45) ) begin
      W_mem_9_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_10_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_48) ) begin
      W_mem_10_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_11_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_49) ) begin
      W_mem_11_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_12_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_50) ) begin
      W_mem_12_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_13_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_51) ) begin
      W_mem_13_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_14_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_52) ) begin
      W_mem_14_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_15_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_53) ) begin
      W_mem_15_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_16_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_55) ) begin
      W_mem_16_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_17_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_57) ) begin
      W_mem_17_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_18_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_58) ) begin
      W_mem_18_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_19_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_59) ) begin
      W_mem_19_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_20_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_61) ) begin
      W_mem_20_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_21_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_63) ) begin
      W_mem_21_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_22_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_64) ) begin
      W_mem_22_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_23_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_65) ) begin
      W_mem_23_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_24_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_66) ) begin
      W_mem_24_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_25_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_67) ) begin
      W_mem_25_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_26_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_68) ) begin
      W_mem_26_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_27_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_69) ) begin
      W_mem_27_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_28_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_70) ) begin
      W_mem_28_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_29_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_71) ) begin
      W_mem_29_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_30_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_72) ) begin
      W_mem_30_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mem_31_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_73) ) begin
      W_mem_31_sva <= W_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mac_pntr_sva <= 5'b00000;
      I_mac_pntr_sva <= 5'b00000;
      O_mac_pntr_sva <= 5'b00000;
      W_irrel_cnt_sva_0 <= 1'b0;
      I_irrel_cnt_sva_0 <= 1'b0;
      O_mac_counter_4_sva <= 5'b00000;
      O_mac_counter_3_sva <= 5'b00000;
      O_mac_counter_2_sva <= 5'b00000;
      O_mac_counter_1_sva <= 5'b00000;
      O_mac_counter_0_sva <= 5'b00000;
      W_mac_counter_4_sva <= 5'b00000;
      W_mac_counter_3_sva <= 5'b00000;
      W_mac_counter_2_sva <= 5'b00000;
      W_mac_counter_1_sva <= 5'b00000;
      W_mac_counter_0_sva <= 5'b00000;
      I_mac_counter_4_sva <= 5'b00000;
      I_mac_counter_3_sva <= 5'b00000;
      I_mac_counter_2_sva <= 5'b00000;
      I_mac_counter_1_sva <= 5'b00000;
      I_mac_counter_0_sva <= 5'b00000;
    end
    else if ( W_mac_pntr_and_cse ) begin
      W_mac_pntr_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_19;
      I_mac_pntr_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_20;
      O_mac_pntr_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_18;
      W_irrel_cnt_sva_0 <= (W_irrel_cnt_sva_dfm_mx0[0]) & if_6_unequal_tmp_2;
      I_irrel_cnt_sva_0 <= (I_irrel_cnt_sva_dfm_mx0[0]) & if_6_unequal_tmp_3;
      O_mac_counter_4_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_24[24:20];
      O_mac_counter_3_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_24[19:15];
      O_mac_counter_2_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_24[14:10];
      O_mac_counter_1_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_24[9:5];
      O_mac_counter_0_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_24[4:0];
      W_mac_counter_4_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_29[24:20];
      W_mac_counter_3_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_29[19:15];
      W_mac_counter_2_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_29[14:10];
      W_mac_counter_1_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_29[9:5];
      W_mac_counter_0_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_29[4:0];
      I_mac_counter_4_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_34[24:20];
      I_mac_counter_3_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_34[19:15];
      I_mac_counter_2_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_34[14:10];
      I_mac_counter_1_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_34[9:5];
      I_mac_counter_0_sva <= libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_34[4:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_0_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_80) ) begin
      I_mem_0_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_1_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_88) ) begin
      I_mem_1_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_2_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_91) ) begin
      I_mem_2_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_3_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_92) ) begin
      I_mem_3_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_4_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_95) ) begin
      I_mem_4_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_5_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_98) ) begin
      I_mem_5_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_6_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_99) ) begin
      I_mem_6_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_7_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_100) ) begin
      I_mem_7_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_8_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_103) ) begin
      I_mem_8_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_9_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_104) ) begin
      I_mem_9_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_10_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_107) ) begin
      I_mem_10_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_11_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_108) ) begin
      I_mem_11_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_12_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_109) ) begin
      I_mem_12_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_13_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_110) ) begin
      I_mem_13_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_14_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_111) ) begin
      I_mem_14_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_15_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_112) ) begin
      I_mem_15_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_16_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_114) ) begin
      I_mem_16_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_17_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_115) ) begin
      I_mem_17_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_18_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_117) ) begin
      I_mem_18_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_19_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_118) ) begin
      I_mem_19_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_20_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_119) ) begin
      I_mem_20_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_21_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_120) ) begin
      I_mem_21_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_22_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_121) ) begin
      I_mem_22_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_23_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_122) ) begin
      I_mem_23_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_24_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_124) ) begin
      I_mem_24_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_25_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_125) ) begin
      I_mem_25_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_26_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_127) ) begin
      I_mem_26_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_27_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_128) ) begin
      I_mem_27_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_28_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_129) ) begin
      I_mem_28_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_29_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_130) ) begin
      I_mem_29_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_30_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_131) ) begin
      I_mem_30_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_mem_31_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_dcpl_132) ) begin
      I_mem_31_sva <= I_wr_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      else_3_land_lpi_1_dfm <= 1'b0;
    end
    else if ( run_wen & (~(mux_419_nl | ((mux_tmp_84 | (~ main_stage_0_2)) & (fsm_output[0]))))
        ) begin
      else_3_land_lpi_1_dfm <= else_3_land_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_0_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_138)) ) begin
      O_mem_0_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_1_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_143)) ) begin
      O_mem_1_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_2_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_147)) ) begin
      O_mem_2_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_3_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_151)) ) begin
      O_mem_3_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_4_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_155)) ) begin
      O_mem_4_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_5_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_158)) ) begin
      O_mem_5_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_6_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_161)) ) begin
      O_mem_6_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_7_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_164)) ) begin
      O_mem_7_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_8_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_168)) ) begin
      O_mem_8_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_9_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_171)) ) begin
      O_mem_9_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_10_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_174)) ) begin
      O_mem_10_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_11_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_177)) ) begin
      O_mem_11_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_12_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_181)) ) begin
      O_mem_12_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_13_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_184)) ) begin
      O_mem_13_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_14_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_187)) ) begin
      O_mem_14_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_15_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_139 | or_dcpl_190)) ) begin
      O_mem_15_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_16_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_138)) ) begin
      O_mem_16_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_17_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_143)) ) begin
      O_mem_17_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_18_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_147)) ) begin
      O_mem_18_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_19_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_151)) ) begin
      O_mem_19_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_20_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_155)) ) begin
      O_mem_20_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_21_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_158)) ) begin
      O_mem_21_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_22_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_161)) ) begin
      O_mem_22_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_23_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_164)) ) begin
      O_mem_23_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_24_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_168)) ) begin
      O_mem_24_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_25_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_171)) ) begin
      O_mem_25_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_26_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_174)) ) begin
      O_mem_26_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_27_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_177)) ) begin
      O_mem_27_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_28_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_181)) ) begin
      O_mem_28_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_29_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_184)) ) begin
      O_mem_29_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_30_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_187)) ) begin
      O_mem_30_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mem_31_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~((~ mux_426_itm) | or_dcpl_193 | or_dcpl_190)) ) begin
      O_mem_31_sva <= mac_data_data_sva_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      skid_buf_top_regs_data_0_0_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_359_cse) ) begin
      skid_buf_top_regs_data_0_0_sva <= mac_data_data_sva_dfm_2_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      skid_buf_top_regs_data_1_0_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_363_cse) ) begin
      skid_buf_top_regs_data_1_0_sva <= mac_data_data_sva_dfm_2_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      skid_buf_top_regs_data_2_0_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ or_367_cse) ) begin
      skid_buf_top_regs_data_2_0_sva <= mac_data_data_sva_dfm_2_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_write_data_data_sva <= 16'b0000000000000000;
    end
    else if ( land_9_lpi_1_dfm_1_1 & run_wen ) begin
      O_write_data_data_sva <= O_write_data_data_sva_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_wr_pntr_sva <= 5'b00000;
    end
    else if ( run_wen & (~(or_dcpl_19 | (~ main_stage_0_2))) ) begin
      W_wr_pntr_sva <= W_wr_pntr_sva_dfm_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_wr_pntr_sva <= 5'b00000;
    end
    else if ( run_wen & (~(or_dcpl_78 | (~ main_stage_0_2))) ) begin
      I_wr_pntr_sva <= I_wr_pntr_sva_dfm_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      skid_buf_top_rd_ptr_sva_0 <= 1'b0;
      skid_buf_top_rd_ptr_sva_1 <= 1'b0;
    end
    else if ( skid_buf_top_rd_ptr_and_cse ) begin
      skid_buf_top_rd_ptr_sva_0 <= skid_buf_top_pop_skid_buf_top_pop_and_4_itm;
      skid_buf_top_rd_ptr_sva_1 <= skid_buf_top_pop_skid_buf_top_pop_and_2_itm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      skid_buf_top_cnt_sva <= 2'b00;
    end
    else if ( mux_597_nl & and_dcpl_34 & (~ (fsm_output[0])) & run_wen ) begin
      skid_buf_top_cnt_sva <= skid_buf_top_cnt_sva_mx1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      skid_buf_top_wr_ptr_sva_0 <= 1'b0;
      skid_buf_top_wr_ptr_sva_1 <= 1'b0;
    end
    else if ( and_370_cse ) begin
      skid_buf_top_wr_ptr_sva_0 <= skid_buf_top_wr_ptr_sva_0_mx0w0;
      skid_buf_top_wr_ptr_sva_1 <= skid_buf_top_wr_ptr_sva_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_irrel_cnt_sva_4_1 <= 4'b0000;
    end
    else if ( mux_601_nl & run_wen & (~ (fsm_output[0])) ) begin
      W_irrel_cnt_sva_4_1 <= W_irrel_cnt_sva_dfm_mx0[4:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_irrel_cnt_sva_4_1 <= 4'b0000;
    end
    else if ( mux_605_nl & run_wen & (~ (fsm_output[0])) ) begin
      I_irrel_cnt_sva_4_1 <= I_irrel_cnt_sva_dfm_mx0[4:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_instr_in_crt_lpi_1_dfm <= 50'b00000000000000000000000000000000000000000000000000;
      I_instr_in_crt_lpi_1_dfm_1 <= 50'b00000000000000000000000000000000000000000000000000;
      W_instr_in_crt_lpi_1_dfm_1 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( and_dcpl_58 ) begin
      O_instr_in_crt_lpi_1_dfm <= O_instr_in_crt_lpi_1_dfm_mx0;
      I_instr_in_crt_lpi_1_dfm_1 <= I_instr_in_crt_lpi_1_dfm_1_mx0;
      W_instr_in_crt_lpi_1_dfm_1 <= W_instr_in_crt_lpi_1_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_vld_zg_pntr_sva <= 5'b00000;
    end
    else if ( mux_614_nl & run_wen & (~ (fsm_output[0])) ) begin
      O_vld_zg_pntr_sva <= if_6_if_6_mux1h_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_data_vld_sva <= 1'b0;
    end
    else if ( run_wen & ((~(and_dcpl_28 | ((~((~((~ mux_460_cse) & or_dcpl_14 & aif_7_equal_tmp))
        & main_stage_0_2)) & (fsm_output[0])))) | O_data_vld_sva_mx0c1) ) begin
      O_data_vld_sva <= MUX_s_1_2_2(O_data_vld_sva_dfm_4_mx0w0, else_8_else_8_or_2_nl,
          O_data_vld_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      else_8_land_lpi_1_dfm <= 1'b0;
    end
    else if ( run_wen & mux_490_nl & (~((~(mux_517_nl & main_stage_0_2)) & (fsm_output[0])))
        ) begin
      else_8_land_lpi_1_dfm <= else_8_land_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_mac_irrel_at_maxBuf_sva <= 1'b0;
      I_mac_irrel_at_maxBuf_sva <= 1'b0;
    end
    else if ( W_mac_irrel_at_maxBuf_and_cse ) begin
      W_mac_irrel_at_maxBuf_sva <= MUX_s_1_2_2(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_26,
          if_for_if_for_and_28_tmp, mux_tmp_76);
      I_mac_irrel_at_maxBuf_sva <= MUX_s_1_2_2(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_31,
          if_for_if_for_and_27_tmp, mux_tmp_76);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mac_tile_bound_4_lpi_1 <= 5'b00000;
      O_mac_tile_bound_3_lpi_1 <= 5'b00000;
      O_mac_tile_bound_2_lpi_1 <= 5'b00000;
      O_mac_tile_bound_1_lpi_1 <= 5'b00000;
      O_mac_tile_bound_0_lpi_1 <= 5'b00000;
      W_mac_tile_bound_4_lpi_1 <= 5'b00000;
      W_mac_tile_bound_3_lpi_1 <= 5'b00000;
      W_mac_tile_bound_2_lpi_1 <= 5'b00000;
      W_mac_tile_bound_1_lpi_1 <= 5'b00000;
      W_mac_tile_bound_0_lpi_1 <= 5'b00000;
      I_mac_tile_bound_4_lpi_1 <= 5'b00000;
      I_mac_tile_bound_3_lpi_1 <= 5'b00000;
      I_mac_tile_bound_2_lpi_1 <= 5'b00000;
      I_mac_tile_bound_1_lpi_1 <= 5'b00000;
      I_mac_tile_bound_0_lpi_1 <= 5'b00000;
    end
    else if ( and_395_cse ) begin
      O_mac_tile_bound_4_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_25[24:20]),
          O_mac_tile_bound_4_lpi_1_dfm_mx0, mux_tmp_76);
      O_mac_tile_bound_3_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_25[19:15]),
          O_mac_tile_bound_3_lpi_1_dfm_mx0, mux_tmp_76);
      O_mac_tile_bound_2_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_25[14:10]),
          O_mac_tile_bound_2_lpi_1_dfm_mx0, mux_tmp_76);
      O_mac_tile_bound_1_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_25[9:5]),
          O_mac_tile_bound_1_lpi_1_dfm_mx0, mux_tmp_76);
      O_mac_tile_bound_0_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_25[4:0]),
          O_mac_tile_bound_0_lpi_1_dfm_mx0, mux_tmp_76);
      W_mac_tile_bound_4_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_30[24:20]),
          W_mac_tile_bound_4_lpi_1_dfm_mx0, mux_tmp_76);
      W_mac_tile_bound_3_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_30[19:15]),
          W_mac_tile_bound_3_lpi_1_dfm_mx0, mux_tmp_76);
      W_mac_tile_bound_2_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_30[14:10]),
          W_mac_tile_bound_2_lpi_1_dfm_mx0, mux_tmp_76);
      W_mac_tile_bound_1_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_30[9:5]),
          W_mac_tile_bound_1_lpi_1_dfm_mx0, mux_tmp_76);
      W_mac_tile_bound_0_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_30[4:0]),
          W_mac_tile_bound_0_lpi_1_dfm_mx0, mux_tmp_76);
      I_mac_tile_bound_4_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_35[24:20]),
          I_mac_tile_bound_4_lpi_1_dfm_mx0, mux_tmp_76);
      I_mac_tile_bound_3_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_35[19:15]),
          I_mac_tile_bound_3_lpi_1_dfm_mx0, mux_tmp_76);
      I_mac_tile_bound_2_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_35[14:10]),
          I_mac_tile_bound_2_lpi_1_dfm_mx0, mux_tmp_76);
      I_mac_tile_bound_1_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_35[9:5]),
          I_mac_tile_bound_1_lpi_1_dfm_mx0, mux_tmp_76);
      I_mac_tile_bound_0_lpi_1 <= MUX_v_5_2_2((libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_35[4:0]),
          I_mac_tile_bound_0_lpi_1_dfm_mx0, mux_tmp_76);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_write_flag_sva <= 1'b0;
    end
    else if ( (~ W_data_vld_sva_dfm_1_1) & run_wen ) begin
      W_write_flag_sva <= W_write_flag_sva_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_write_flag_sva <= 1'b0;
    end
    else if ( (~ I_data_vld_sva_dfm_1_1) & run_wen ) begin
      I_write_flag_sva <= I_write_flag_sva_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      skid_buf_top_cnt_sva_1_1 <= 2'b00;
      skid_buf_top_wr_ptr_sva_dfm_1_1 <= 1'b0;
    end
    else if ( skid_buf_top_cnt_and_1_cse ) begin
      skid_buf_top_cnt_sva_1_1 <= nl_skid_buf_top_cnt_sva_1_1[1:0];
      skid_buf_top_wr_ptr_sva_dfm_1_1 <= skid_buf_top_push_and_psp_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      if_5_if_nbw_stat_sva <= 1'b0;
    end
    else if ( flags_wr_zero_guard_and_cse & ((~ mux_341_nl) | (~ O_mac_irrel_at_max_sva_dfm_mx0)
        | flags_top_1_1_sva) & (~(or_dcpl_226 | (~ if_5_and_svs_1))) ) begin
      if_5_if_nbw_stat_sva <= O_rd_data_rsci_irdy_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      I_vld_pntr_sva_dfm_1_1 <= 5'b00000;
    end
    else if ( run_wen & (~(main_stage_0_2 & (~ mux_530_itm))) ) begin
      I_vld_pntr_sva_dfm_1_1 <= MUX_v_5_2_2(5'b00000, libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_20,
          mux_530_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      W_vld_pntr_sva_dfm_1_1 <= 5'b00000;
    end
    else if ( run_wen & (~(main_stage_0_2 & (~ mux_543_itm))) ) begin
      W_vld_pntr_sva_dfm_1_1 <= MUX_v_5_2_2(5'b00000, libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_19,
          mux_543_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      aif_2_land_1_lpi_1_dfm <= 1'b0;
      aif_3_land_lpi_1_dfm <= 1'b0;
    end
    else if ( and_426_cse ) begin
      aif_2_land_1_lpi_1_dfm <= aif_2_land_1_lpi_1_dfm_mx0;
      aif_3_land_lpi_1_dfm <= aif_3_land_lpi_1_dfm_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      O_mac_irrel_at_max_sva <= 1'b1;
    end
    else if ( mux_672_nl & run_wen ) begin
      O_mac_irrel_at_max_sva <= MUX_s_1_2_2(libraries_O_addr_cnt_5_O_addr_type_L1_1_7448a59bcc55848f49259c21df88d8bc12ff1_21,
          O_mac_irrel_at_max_sva_dfm_mx0, or_531_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      skid_buf_wr_zero_guard_regs_1_sva_dfm_1 <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_246) ) begin
      skid_buf_wr_zero_guard_regs_1_sva_dfm_1 <= wr_data_zero_guard_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      skid_buf_wr_zero_guard_regs_0_sva_dfm_1 <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_248 | (fsm_output[0]))) ) begin
      skid_buf_wr_zero_guard_regs_0_sva_dfm_1 <= wr_data_zero_guard_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      skid_buf_wr_zero_guard_cnt_sva <= 2'b00;
    end
    else if ( (mux_675_nl | and_432_cse) & (~ (fsm_output[0])) & run_wen ) begin
      skid_buf_wr_zero_guard_cnt_sva <= mux1h_1_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      skid_buf_wr_zero_guard_wr_ptr_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_tmp_162 | (fsm_output[0]))) ) begin
      skid_buf_wr_zero_guard_wr_ptr_sva <= ~ skid_buf_wr_zero_guard_wr_ptr_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      skid_buf_wr_zero_guard_rd_ptr_sva <= 1'b0;
    end
    else if ( run_wen & ((else_8_land_lpi_1_dfm_mx0w0 & (~ (fsm_output[0]))) | or_tmp_242)
        ) begin
      skid_buf_wr_zero_guard_rd_ptr_sva <= ~ skid_buf_wr_zero_guard_rd_ptr_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      flags_top_1_1_sva <= 1'b0;
    end
    else if ( run_wen & (main_stage_0_2 | flags_top_1_1_sva_mx0c1) ) begin
      flags_top_1_1_sva <= ~((~((mux1h_7_tmp!=2'b00))) | flags_top_1_1_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      skid_buf_top_push_nor_psp <= 1'b0;
      skid_buf_top_push_and_psp <= 1'b0;
      skid_buf_top_push_and_1_psp <= 1'b0;
    end
    else if ( skid_buf_top_push_and_2_cse ) begin
      skid_buf_top_push_nor_psp <= skid_buf_top_push_nor_psp_mx0w0;
      skid_buf_top_push_and_psp <= skid_buf_top_push_and_psp_1;
      skid_buf_top_push_and_1_psp <= skid_buf_top_push_and_1_psp_mx0w0;
    end
  end
  assign nor_182_nl = ~(and_526_cse | (W_irrel_cnt_sva_4_1!=4'b0000) | not_tmp_9);
  assign nor_183_nl = ~(and_526_cse | (if_6_if_3_acc_tmp[4:1]!=4'b0000) | not_tmp_8);
  assign mux_354_nl = MUX_s_1_2_2(nor_182_nl, nor_183_nl, W_mac_irrel_at_maxBuf_sva);
  assign nor_184_nl = ~(nor_tmp_8 | (W_irrel_cnt_sva_4_1!=4'b0000) | not_tmp_9);
  assign nor_185_nl = ~(nor_tmp_8 | (if_6_if_3_acc_tmp[4:1]!=4'b0000) | not_tmp_8);
  assign mux_353_nl = MUX_s_1_2_2(nor_184_nl, nor_185_nl, if_for_if_for_and_28_tmp);
  assign mux_355_nl = MUX_s_1_2_2(mux_354_nl, mux_353_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign nor_178_nl = ~(and_526_cse | (I_irrel_cnt_sva_4_1!=4'b0000) | not_tmp_15);
  assign nor_179_nl = ~(and_526_cse | (if_6_if_1_acc_tmp[4:1]!=4'b0000) | not_tmp_14);
  assign mux_359_nl = MUX_s_1_2_2(nor_178_nl, nor_179_nl, I_mac_irrel_at_maxBuf_sva);
  assign nor_180_nl = ~(nor_tmp_8 | (I_irrel_cnt_sva_4_1!=4'b0000) | not_tmp_15);
  assign nor_181_nl = ~(nor_tmp_8 | (if_6_if_1_acc_tmp[4:1]!=4'b0000) | not_tmp_14);
  assign mux_358_nl = MUX_s_1_2_2(nor_180_nl, nor_181_nl, if_for_if_for_and_27_tmp);
  assign mux_360_nl = MUX_s_1_2_2(mux_359_nl, mux_358_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign mux_386_nl = MUX_s_1_2_2(or_18_cse, or_tmp_73, nor_tmp_26);
  assign mux_385_nl = MUX_s_1_2_2(or_18_cse, or_tmp_73, nor_tmp_25);
  assign mux_387_nl = MUX_s_1_2_2(mux_386_nl, mux_385_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign and_293_nl = O_mac_irrel_at_max_sva & and_306_cse;
  assign and_294_nl = if_for_if_for_and_26_tmp & and_306_cse;
  assign mux_384_nl = MUX_s_1_2_2(and_293_nl, and_294_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign or_97_nl = (mux1h_7_tmp!=2'b00) | mux_384_nl;
  assign mux_388_nl = MUX_s_1_2_2(mux_387_nl, or_97_nl, main_stage_0_2);
  assign if_6_if_6_and_3_nl = W_data_vld_sva_mx0 & if_6_unequal_tmp_2;
  assign if_6_if_6_and_nl = I_data_vld_sva_mx0 & if_6_unequal_tmp_3;
  assign if_6_if_6_and_9_nl = O_write_flag_sva_mx0 & land_lpi_1_dfm_1;
  assign if_6_if_if_6_if_and_nl = data_zg_sva & (~ if_6_else_if_equal_tmp);
  assign if_6_mux_3_nl = MUX_s_1_2_2(data_zg_sva, if_6_if_if_6_if_and_nl, land_lpi_1_dfm_1);
  assign mux_123_nl = MUX_s_1_2_2(data_zg_sva, if_6_mux_3_nl, lor_4_lpi_1_dfm_1);
  assign if_5_if_or_nl = ((((~ or_360_tmp) & skid_buf_top_peek_and_m1c) | ((~ or_364_tmp)
      & skid_buf_top_peek_and_4_m1c) | ((~ or_368_tmp) & skid_buf_top_peek_and_5_m1c))
      & O_rd_data_rsci_idat_mx0c0) | ((~ or_359_cse) & if_5_if_and_3_m1c) | ((~ or_363_cse)
      & if_5_if_and_4_m1c) | ((~ or_367_cse) & if_5_if_and_5_m1c);
  assign if_5_if_or_2_nl = (or_360_tmp & skid_buf_top_peek_and_m1c & O_rd_data_rsci_idat_mx0c0)
      | (or_359_cse & if_5_if_and_3_m1c);
  assign if_5_if_or_3_nl = (((skid_buf_top_push_nor_psp_mx0w0 & skid_buf_top_peek_nor_m1c_1)
      | (skid_buf_top_push_and_psp_1 & skid_buf_top_peek_and_m1c_2) | (skid_buf_top_push_and_1_psp_mx0w0
      & skid_buf_top_peek_and_m1c_3)) & O_rd_data_rsci_idat_mx0c0) | O_rd_data_rsci_idat_mx0c2;
  assign if_5_if_or_4_nl = (or_364_tmp & skid_buf_top_peek_and_4_m1c & O_rd_data_rsci_idat_mx0c0)
      | (or_363_cse & if_5_if_and_4_m1c);
  assign if_5_if_or_5_nl = (or_368_tmp & skid_buf_top_peek_and_5_m1c & O_rd_data_rsci_idat_mx0c0)
      | (or_367_cse & if_5_if_and_5_m1c);
  assign nand_37_nl = ~(oif_1_unequal_tmp & oif_2_unequal_tmp & oif_unequal_tmp &
      (~ and_tmp_56));
  assign nand_36_nl = ~(oif_1_unequal_tmp & oif_2_unequal_tmp & (~ and_tmp_56));
  assign mux_418_nl = MUX_s_1_2_2(nand_37_nl, nand_36_nl, O_data_vld_sva);
  assign nor_175_nl = ~(land_lpi_1_dfm_1 | mux_418_nl);
  assign mux_419_nl = MUX_s_1_2_2(nor_175_nl, mux_tmp_84, main_stage_0_2);
  assign mux_595_nl = MUX_s_1_2_2(or_tmp_299, mux_tmp_251, and_541_cse);
  assign mux_596_nl = MUX_s_1_2_2(mux_595_nl, mux_tmp_251, or_tmp_300);
  assign or_593_nl = (~ O_mac_irrel_at_max_sva) | flags_top_1_1_sva;
  assign mux_597_nl = MUX_s_1_2_2(mux_596_nl, or_tmp_299, or_593_nl);
  assign and_537_nl = oif_2_unequal_tmp & or_1_cse & oif_1_unequal_tmp & not_tmp_165;
  assign nand_101_nl = ~(mux_124_itm_1 & (~ nand_tmp_39));
  assign nand_100_nl = ~(O_wr_data_rsci_ivld_mxwt & (~ nand_tmp_39));
  assign mux_599_nl = MUX_s_1_2_2(nand_101_nl, nand_100_nl, land_9_lpi_1_dfm_1_1);
  assign mux_600_nl = MUX_s_1_2_2(mux_599_nl, nand_tmp_39, or_1_cse);
  assign nor_302_nl = ~(nor_303_cse | mux_600_nl);
  assign mux_601_nl = MUX_s_1_2_2(and_537_nl, nor_302_nl, main_stage_0_2);
  assign and_533_nl = oif_2_unequal_tmp & or_1_cse & oif_1_unequal_tmp & not_tmp_172;
  assign nand_108_nl = ~(mux_124_itm_1 & (~ nand_tmp_46));
  assign nand_107_nl = ~(O_wr_data_rsci_ivld_mxwt & (~ nand_tmp_46));
  assign mux_603_nl = MUX_s_1_2_2(nand_108_nl, nand_107_nl, land_9_lpi_1_dfm_1_1);
  assign mux_604_nl = MUX_s_1_2_2(mux_603_nl, nand_tmp_46, or_1_cse);
  assign nor_299_nl = ~(nor_303_cse | mux_604_nl);
  assign mux_605_nl = MUX_s_1_2_2(and_533_nl, nor_299_nl, main_stage_0_2);
  assign and_388_nl = oif_2_unequal_tmp & oif_1_unequal_tmp & nor_tmp_189;
  assign mux_611_nl = MUX_s_1_2_2(and_tmp_107, or_tmp_10, mux_124_itm_1);
  assign mux_610_nl = MUX_s_1_2_2(and_tmp_107, or_tmp_10, O_wr_data_rsci_ivld_mxwt);
  assign mux_612_nl = MUX_s_1_2_2(mux_611_nl, mux_610_nl, land_9_lpi_1_dfm_1_1);
  assign and_387_nl = or_620_cse & mux_612_nl;
  assign mux_613_nl = MUX_s_1_2_2(and_388_nl, and_387_nl, main_stage_0_2);
  assign and_385_nl = oif_2_unequal_tmp & oif_1_unequal_tmp & and_tmp_103;
  assign mux_607_nl = MUX_s_1_2_2(and_tmp_104, and_tmp_102, mux_124_itm_1);
  assign mux_606_nl = MUX_s_1_2_2(and_tmp_104, and_tmp_102, O_wr_data_rsci_ivld_mxwt);
  assign mux_608_nl = MUX_s_1_2_2(mux_607_nl, mux_606_nl, land_9_lpi_1_dfm_1_1);
  assign and_384_nl = or_620_cse & mux_608_nl;
  assign mux_609_nl = MUX_s_1_2_2(and_385_nl, and_384_nl, main_stage_0_2);
  assign mux_614_nl = MUX_s_1_2_2(mux_613_nl, mux_609_nl, and_526_cse);
  assign else_8_else_8_or_2_nl = O_data_vld_sva_dfm_4_mx0 | else_8_land_lpi_1_dfm_mx0w0;
  assign mux_488_nl = MUX_s_1_2_2(mux_tmp_153, mux_tmp_143, mux_124_itm_1);
  assign mux_487_nl = MUX_s_1_2_2(mux_tmp_153, mux_tmp_143, O_wr_data_rsci_ivld_mxwt);
  assign mux_489_nl = MUX_s_1_2_2(mux_488_nl, mux_487_nl, land_9_lpi_1_dfm_1_1);
  assign mux_490_nl = MUX_s_1_2_2(mux_tmp_153, mux_489_nl, nor_108_cse);
  assign mux_515_nl = MUX_s_1_2_2(mux_tmp_180, mux_tmp_170, mux_124_itm_1);
  assign mux_514_nl = MUX_s_1_2_2(mux_tmp_180, mux_tmp_170, O_wr_data_rsci_ivld_mxwt);
  assign mux_516_nl = MUX_s_1_2_2(mux_515_nl, mux_514_nl, land_9_lpi_1_dfm_1_1);
  assign mux_517_nl = MUX_s_1_2_2(mux_tmp_180, mux_516_nl, nor_108_cse);
  assign nl_skid_buf_top_cnt_sva_1_1  = skid_buf_top_cnt_sva_mx1 + 2'b01;
  assign and_52_nl = or_558_cse & mux_tmp_6;
  assign mux_340_nl = MUX_s_1_2_2(and_52_nl, mux_tmp_6, oif_2_unequal_tmp);
  assign and_49_nl = or_558_cse & mux_tmp_4;
  assign mux_335_nl = MUX_s_1_2_2(and_tmp_1, and_tmp, I_data_vld_sva_dfm_1_1);
  assign mux_336_nl = MUX_s_1_2_2(mux_335_nl, mux_554_cse, oif_1_unequal_tmp);
  assign mux_338_nl = MUX_s_1_2_2(and_49_nl, mux_336_nl, oif_2_unequal_tmp);
  assign mux_341_nl = MUX_s_1_2_2(mux_340_nl, mux_338_nl, or_1_cse);
  assign or_555_nl = and_526_cse | (~ mux_tmp_14);
  assign or_556_nl = nor_tmp_8 | (~ mux_tmp_14);
  assign mux_553_nl = MUX_s_1_2_2(or_555_nl, or_556_nl, reg_W_instr_in_rsci_oswt_cse_1);
  assign or_531_nl = (mux_tmp_76 & (fsm_output[1])) | (mux_553_nl & main_stage_0_2);
  assign mux_716_nl = MUX_s_1_2_2((fsm_output[1]), nor_tmp_217, and_526_cse);
  assign mux_670_nl = MUX_s_1_2_2(nor_tmp_217, mux_716_nl, and_544_cse);
  assign mux_671_nl = MUX_s_1_2_2(nor_tmp_217, mux_670_nl, oif_2_unequal_tmp);
  assign mux_721_nl = MUX_s_1_2_2(reg_W_instr_in_rsci_oswt_cse_1, mux_663_itm, or_tmp_10);
  assign mux_666_nl = MUX_s_1_2_2(reg_W_instr_in_rsci_oswt_cse_1, mux_721_nl, mux_124_itm_1);
  assign mux_722_nl = MUX_s_1_2_2(reg_W_instr_in_rsci_oswt_cse_1, mux_663_itm, or_tmp_10);
  assign mux_665_nl = MUX_s_1_2_2(reg_W_instr_in_rsci_oswt_cse_1, mux_722_nl, O_wr_data_rsci_ivld_mxwt);
  assign mux_667_nl = MUX_s_1_2_2(mux_666_nl, mux_665_nl, land_9_lpi_1_dfm_1_1);
  assign mux_664_nl = MUX_s_1_2_2(reg_W_instr_in_rsci_oswt_cse_1, mux_663_itm, or_tmp_10);
  assign mux_668_nl = MUX_s_1_2_2(mux_667_nl, mux_664_nl, or_1_cse);
  assign mux_669_nl = MUX_s_1_2_2(reg_W_instr_in_rsci_oswt_cse_1, mux_668_nl, or_620_cse);
  assign mux_672_nl = MUX_s_1_2_2(mux_671_nl, mux_669_nl, main_stage_0_2);
  assign or_757_nl = (~(mux_404_tmp | (~(else_8_land_lpi_1_dfm & ((skid_buf_wr_zero_guard_cnt_sva!=2'b00))))))
      | land_8_lpi_1_dfm_1;
  assign mux_675_nl = MUX_s_1_2_2(land_8_lpi_1_dfm_1, or_757_nl, aif_7_equal_tmp);
  assign UPDATE_PSUM_FROM_TOP_or_2_nl = (~((~(or_dcpl_25 | or_dcpl_23)) | and_331_cse))
      | (or_dcpl_21 & and_331_cse);
  assign UPDATE_PSUM_FROM_TOP_mux_5_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_0_sva,
      UPDATE_PSUM_FROM_TOP_or_2_nl);
  assign if_10_mux_97_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_1_sva, or_dcpl_29);
  assign if_10_mux_98_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_2_sva, or_dcpl_32);
  assign if_10_mux_99_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_3_sva, or_dcpl_33);
  assign if_10_mux_100_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_4_sva, or_dcpl_36);
  assign if_10_mux_101_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_5_sva, or_dcpl_39);
  assign if_10_mux_102_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_6_sva, or_dcpl_40);
  assign if_10_mux_103_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_7_sva, or_dcpl_41);
  assign if_10_mux_104_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_8_sva, or_dcpl_44);
  assign if_10_mux_105_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_9_sva, or_dcpl_45);
  assign if_10_mux_106_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_10_sva,
      or_dcpl_48);
  assign if_10_mux_107_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_11_sva,
      or_dcpl_49);
  assign if_10_mux_108_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_12_sva,
      or_dcpl_50);
  assign if_10_mux_109_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_13_sva,
      or_dcpl_51);
  assign if_10_mux_110_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_14_sva,
      or_dcpl_52);
  assign if_10_mux_111_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_15_sva,
      or_dcpl_53);
  assign if_10_mux_112_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_16_sva,
      or_dcpl_55);
  assign if_10_mux_113_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_17_sva,
      or_dcpl_57);
  assign if_10_mux_114_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_18_sva,
      or_dcpl_58);
  assign if_10_mux_115_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_19_sva,
      or_dcpl_59);
  assign if_10_mux_116_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_20_sva,
      or_dcpl_61);
  assign if_10_mux_117_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_21_sva,
      or_dcpl_63);
  assign if_10_mux_118_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_22_sva,
      or_dcpl_64);
  assign if_10_mux_119_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_23_sva,
      or_dcpl_65);
  assign if_10_mux_120_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_24_sva,
      or_dcpl_66);
  assign if_10_mux_121_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_25_sva,
      or_dcpl_67);
  assign if_10_mux_122_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_26_sva,
      or_dcpl_68);
  assign if_10_mux_123_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_27_sva,
      or_dcpl_69);
  assign if_10_mux_124_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_28_sva,
      or_dcpl_70);
  assign if_10_mux_125_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_29_sva,
      or_dcpl_71);
  assign if_10_mux_126_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_30_sva,
      or_dcpl_72);
  assign if_10_mux_127_nl = MUX_v_16_2_2(W_wr_data_rsci_idat_mxwt, W_mem_31_sva,
      or_dcpl_73);
  assign mux_723_nl = MUX_v_16_32_2(UPDATE_PSUM_FROM_TOP_mux_5_nl, if_10_mux_97_nl,
      if_10_mux_98_nl, if_10_mux_99_nl, if_10_mux_100_nl, if_10_mux_101_nl, if_10_mux_102_nl,
      if_10_mux_103_nl, if_10_mux_104_nl, if_10_mux_105_nl, if_10_mux_106_nl, if_10_mux_107_nl,
      if_10_mux_108_nl, if_10_mux_109_nl, if_10_mux_110_nl, if_10_mux_111_nl, if_10_mux_112_nl,
      if_10_mux_113_nl, if_10_mux_114_nl, if_10_mux_115_nl, if_10_mux_116_nl, if_10_mux_117_nl,
      if_10_mux_118_nl, if_10_mux_119_nl, if_10_mux_120_nl, if_10_mux_121_nl, if_10_mux_122_nl,
      if_10_mux_123_nl, if_10_mux_124_nl, if_10_mux_125_nl, if_10_mux_126_nl, if_10_mux_127_nl,
      W_mac_pntr_sva);
  assign UPDATE_PSUM_FROM_TOP_or_3_nl = (~((~(or_dcpl_84 | or_dcpl_82)) | and_331_cse))
      | (or_dcpl_80 & and_331_cse);
  assign UPDATE_PSUM_FROM_TOP_mux_6_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_0_sva,
      UPDATE_PSUM_FROM_TOP_or_3_nl);
  assign if_9_mux_97_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_1_sva, or_dcpl_88);
  assign if_9_mux_98_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_2_sva, or_dcpl_91);
  assign if_9_mux_99_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_3_sva, or_dcpl_92);
  assign if_9_mux_100_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_4_sva, or_dcpl_95);
  assign if_9_mux_101_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_5_sva, or_dcpl_98);
  assign if_9_mux_102_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_6_sva, or_dcpl_99);
  assign if_9_mux_103_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_7_sva, or_dcpl_100);
  assign if_9_mux_104_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_8_sva, or_dcpl_103);
  assign if_9_mux_105_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_9_sva, or_dcpl_104);
  assign if_9_mux_106_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_10_sva, or_dcpl_107);
  assign if_9_mux_107_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_11_sva, or_dcpl_108);
  assign if_9_mux_108_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_12_sva, or_dcpl_109);
  assign if_9_mux_109_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_13_sva, or_dcpl_110);
  assign if_9_mux_110_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_14_sva, or_dcpl_111);
  assign if_9_mux_111_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_15_sva, or_dcpl_112);
  assign if_9_mux_112_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_16_sva, or_dcpl_114);
  assign if_9_mux_113_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_17_sva, or_dcpl_115);
  assign if_9_mux_114_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_18_sva, or_dcpl_117);
  assign if_9_mux_115_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_19_sva, or_dcpl_118);
  assign if_9_mux_116_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_20_sva, or_dcpl_119);
  assign if_9_mux_117_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_21_sva, or_dcpl_120);
  assign if_9_mux_118_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_22_sva, or_dcpl_121);
  assign if_9_mux_119_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_23_sva, or_dcpl_122);
  assign if_9_mux_120_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_24_sva, or_dcpl_124);
  assign if_9_mux_121_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_25_sva, or_dcpl_125);
  assign if_9_mux_122_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_26_sva, or_dcpl_127);
  assign if_9_mux_123_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_27_sva, or_dcpl_128);
  assign if_9_mux_124_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_28_sva, or_dcpl_129);
  assign if_9_mux_125_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_29_sva, or_dcpl_130);
  assign if_9_mux_126_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_30_sva, or_dcpl_131);
  assign if_9_mux_127_nl = MUX_v_16_2_2(I_wr_data_rsci_idat_mxwt, I_mem_31_sva, or_dcpl_132);
  assign mux_724_nl = MUX_v_16_32_2(UPDATE_PSUM_FROM_TOP_mux_6_nl, if_9_mux_97_nl,
      if_9_mux_98_nl, if_9_mux_99_nl, if_9_mux_100_nl, if_9_mux_101_nl, if_9_mux_102_nl,
      if_9_mux_103_nl, if_9_mux_104_nl, if_9_mux_105_nl, if_9_mux_106_nl, if_9_mux_107_nl,
      if_9_mux_108_nl, if_9_mux_109_nl, if_9_mux_110_nl, if_9_mux_111_nl, if_9_mux_112_nl,
      if_9_mux_113_nl, if_9_mux_114_nl, if_9_mux_115_nl, if_9_mux_116_nl, if_9_mux_117_nl,
      if_9_mux_118_nl, if_9_mux_119_nl, if_9_mux_120_nl, if_9_mux_121_nl, if_9_mux_122_nl,
      if_9_mux_123_nl, if_9_mux_124_nl, if_9_mux_125_nl, if_9_mux_126_nl, if_9_mux_127_nl,
      I_mac_pntr_sva);
  assign nl_z_out_2 = mux_723_nl * mux_724_nl;
  assign z_out_2 = nl_z_out_2[15:0];
  assign and_549_nl = if_5_and_svs_1 & (fsm_output[1]);
  assign skid_buf_top_pop_1_mux_1_nl = MUX_v_2_2_2(skid_buf_top_cnt_sva, skid_buf_top_cnt_sva_1_1,
      and_549_nl);
  assign nl_z_out_3 = skid_buf_top_pop_1_mux_1_nl + 2'b11;
  assign z_out_3 = nl_z_out_3[1:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_5_2;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [4:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    result = result | ( input_4 & {16{sel[4]}});
    MUX1HOT_v_16_5_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_32_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [15:0] input_22;
    input [15:0] input_23;
    input [15:0] input_24;
    input [15:0] input_25;
    input [15:0] input_26;
    input [15:0] input_27;
    input [15:0] input_28;
    input [15:0] input_29;
    input [15:0] input_30;
    input [15:0] input_31;
    input [4:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_16_32_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [49:0] MUX_v_50_2_2;
    input [49:0] input_0;
    input [49:0] input_1;
    input [0:0] sel;
    reg [49:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_50_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3
// ------------------------------------------------------------------


module config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3
    (
  clk, rst, layer_instruction_in_rsc_dat, layer_instruction_in_rsc_vld, layer_instruction_in_rsc_rdy,
      O_instr_L1_out_rsc_dat, O_instr_L1_out_rsc_vld, O_instr_L1_out_rsc_rdy, O_instr_L2_out_rsc_dat,
      O_instr_L2_out_rsc_vld, O_instr_L2_out_rsc_rdy, O_instr_L3_out_rsc_dat, O_instr_L3_out_rsc_vld,
      O_instr_L3_out_rsc_rdy, I_instr_L1_out_rsc_dat, I_instr_L1_out_rsc_vld, I_instr_L1_out_rsc_rdy,
      I_instr_L2_out_rsc_dat, I_instr_L2_out_rsc_vld, I_instr_L2_out_rsc_rdy, I_instr_L3_out_rsc_dat,
      I_instr_L3_out_rsc_vld, I_instr_L3_out_rsc_rdy, W_instr_L1_out_rsc_dat, W_instr_L1_out_rsc_vld,
      W_instr_L1_out_rsc_rdy, W_instr_L2_out_rsc_dat, W_instr_L2_out_rsc_vld, W_instr_L2_out_rsc_rdy,
      W_instr_L3_out_rsc_dat, W_instr_L3_out_rsc_vld, W_instr_L3_out_rsc_rdy
);
  input clk;
  input rst;
  input [484:0] layer_instruction_in_rsc_dat;
  input layer_instruction_in_rsc_vld;
  output layer_instruction_in_rsc_rdy;
  output [49:0] O_instr_L1_out_rsc_dat;
  output O_instr_L1_out_rsc_vld;
  input O_instr_L1_out_rsc_rdy;
  output [89:0] O_instr_L2_out_rsc_dat;
  output O_instr_L2_out_rsc_vld;
  input O_instr_L2_out_rsc_rdy;
  output [139:0] O_instr_L3_out_rsc_dat;
  output O_instr_L3_out_rsc_vld;
  input O_instr_L3_out_rsc_rdy;
  output [49:0] I_instr_L1_out_rsc_dat;
  output I_instr_L1_out_rsc_vld;
  input I_instr_L1_out_rsc_rdy;
  output [89:0] I_instr_L2_out_rsc_dat;
  output I_instr_L2_out_rsc_vld;
  input I_instr_L2_out_rsc_rdy;
  output [139:0] I_instr_L3_out_rsc_dat;
  output I_instr_L3_out_rsc_vld;
  input I_instr_L3_out_rsc_rdy;
  output [49:0] W_instr_L1_out_rsc_dat;
  output W_instr_L1_out_rsc_vld;
  input W_instr_L1_out_rsc_rdy;
  output [109:0] W_instr_L2_out_rsc_dat;
  output W_instr_L2_out_rsc_vld;
  input W_instr_L2_out_rsc_rdy;
  output [159:0] W_instr_L3_out_rsc_dat;
  output W_instr_L3_out_rsc_vld;
  input W_instr_L3_out_rsc_rdy;


  // Interconnect Declarations
  wire [79:0] W_tiling_unit_L3_run_cmp_loops_bound_rsc_dat;
  wire [4:0] W_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat;
  wire [15:0] W_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat;
  wire [15:0] W_tiling_unit_L3_run_cmp_tile_size_out_rsc_z;
  wire [79:0] W_tiling_unit_L3_run_cmp_instr_bound_rsc_z;
  wire [79:0] W_tiling_unit_L3_run_cmp_instr_tile_rsc_z;
  wire W_tiling_unit_L3_run_cmp_ccs_ccore_start_rsc_dat;
  wire W_tiling_unit_L3_run_cmp_ccs_ccore_en;
  wire CGHpart_irsig_1;
  wire [54:0] W_tiling_unit_L2_run_cmp_loops_bound_rsc_dat;
  wire [4:0] W_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat;
  wire [10:0] W_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat;
  wire [10:0] W_tiling_unit_L2_run_cmp_tile_size_out_rsc_z;
  wire [54:0] W_tiling_unit_L2_run_cmp_instr_bound_rsc_z;
  wire [54:0] W_tiling_unit_L2_run_cmp_instr_tile_rsc_z;
  wire W_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat;
  wire W_tiling_unit_L2_run_cmp_ccs_ccore_en;
  wire [69:0] O_tiling_unit_L3_run_cmp_loops_bound_rsc_dat;
  wire [4:0] O_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat;
  wire [13:0] O_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat;
  wire [13:0] O_tiling_unit_L3_run_cmp_tile_size_out_rsc_z;
  wire [69:0] O_tiling_unit_L3_run_cmp_instr_bound_rsc_z;
  wire [69:0] O_tiling_unit_L3_run_cmp_instr_tile_rsc_z;
  wire O_tiling_unit_L3_run_cmp_ccs_ccore_en;
  wire [44:0] O_tiling_unit_L2_run_cmp_loops_bound_rsc_dat;
  wire [4:0] O_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat;
  wire [8:0] O_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat;
  wire [8:0] O_tiling_unit_L2_run_cmp_tile_size_out_rsc_z;
  wire [44:0] O_tiling_unit_L2_run_cmp_instr_bound_rsc_z;
  wire [44:0] O_tiling_unit_L2_run_cmp_instr_tile_rsc_z;
  wire O_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat;
  wire O_tiling_unit_L2_run_cmp_ccs_ccore_en;
  wire [24:0] O_tiling_unit_L1_run_cmp_loops_bound_rsc_dat;
  wire [4:0] O_tiling_unit_L1_run_cmp_loops_relevancy_rsc_dat;
  wire [4:0] O_tiling_unit_L1_run_cmp_tile_size_in_rsc_dat;
  wire [4:0] O_tiling_unit_L1_run_cmp_tile_size_out_rsc_z;
  wire [24:0] O_tiling_unit_L1_run_cmp_instr_bound_rsc_z;
  wire [24:0] O_tiling_unit_L1_run_cmp_instr_tile_rsc_z;
  wire O_tiling_unit_L1_run_cmp_ccs_ccore_start_rsc_dat;
  wire O_tiling_unit_L1_run_cmp_ccs_ccore_en;


  // Interconnect Declarations for Component Instantiations 
  tiling_unit_5_W_addr_type_L3  W_tiling_unit_L3_run_cmp (
      .loops_bound_rsc_dat(W_tiling_unit_L3_run_cmp_loops_bound_rsc_dat),
      .loops_relevancy_rsc_dat(W_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat),
      .tile_size_in_rsc_dat(W_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat),
      .tile_size_out_rsc_z(W_tiling_unit_L3_run_cmp_tile_size_out_rsc_z),
      .instr_bound_rsc_z(W_tiling_unit_L3_run_cmp_instr_bound_rsc_z),
      .instr_tile_rsc_z(W_tiling_unit_L3_run_cmp_instr_tile_rsc_z),
      .ccs_ccore_start_rsc_dat(W_tiling_unit_L3_run_cmp_ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(clk),
      .ccs_ccore_srst(rst),
      .ccs_ccore_en(W_tiling_unit_L3_run_cmp_ccs_ccore_en)
    );
  tiling_unit_5_W_addr_type_L2  W_tiling_unit_L2_run_cmp (
      .loops_bound_rsc_dat(W_tiling_unit_L2_run_cmp_loops_bound_rsc_dat),
      .loops_relevancy_rsc_dat(W_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat),
      .tile_size_in_rsc_dat(W_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat),
      .tile_size_out_rsc_z(W_tiling_unit_L2_run_cmp_tile_size_out_rsc_z),
      .instr_bound_rsc_z(W_tiling_unit_L2_run_cmp_instr_bound_rsc_z),
      .instr_tile_rsc_z(W_tiling_unit_L2_run_cmp_instr_tile_rsc_z),
      .ccs_ccore_start_rsc_dat(W_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(clk),
      .ccs_ccore_srst(rst),
      .ccs_ccore_en(W_tiling_unit_L2_run_cmp_ccs_ccore_en)
    );
  tiling_unit_5_O_addr_type_L3  O_tiling_unit_L3_run_cmp (
      .loops_bound_rsc_dat(O_tiling_unit_L3_run_cmp_loops_bound_rsc_dat),
      .loops_relevancy_rsc_dat(O_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat),
      .tile_size_in_rsc_dat(O_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat),
      .tile_size_out_rsc_z(O_tiling_unit_L3_run_cmp_tile_size_out_rsc_z),
      .instr_bound_rsc_z(O_tiling_unit_L3_run_cmp_instr_bound_rsc_z),
      .instr_tile_rsc_z(O_tiling_unit_L3_run_cmp_instr_tile_rsc_z),
      .ccs_ccore_start_rsc_dat(CGHpart_irsig_1),
      .ccs_ccore_clk(clk),
      .ccs_ccore_srst(rst),
      .ccs_ccore_en(O_tiling_unit_L3_run_cmp_ccs_ccore_en)
    );
  tiling_unit_5_O_addr_type_L2  O_tiling_unit_L2_run_cmp (
      .loops_bound_rsc_dat(O_tiling_unit_L2_run_cmp_loops_bound_rsc_dat),
      .loops_relevancy_rsc_dat(O_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat),
      .tile_size_in_rsc_dat(O_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat),
      .tile_size_out_rsc_z(O_tiling_unit_L2_run_cmp_tile_size_out_rsc_z),
      .instr_bound_rsc_z(O_tiling_unit_L2_run_cmp_instr_bound_rsc_z),
      .instr_tile_rsc_z(O_tiling_unit_L2_run_cmp_instr_tile_rsc_z),
      .ccs_ccore_start_rsc_dat(O_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(clk),
      .ccs_ccore_srst(rst),
      .ccs_ccore_en(O_tiling_unit_L2_run_cmp_ccs_ccore_en)
    );
  tiling_unit_5_O_addr_type_L1  O_tiling_unit_L1_run_cmp (
      .loops_bound_rsc_dat(O_tiling_unit_L1_run_cmp_loops_bound_rsc_dat),
      .loops_relevancy_rsc_dat(O_tiling_unit_L1_run_cmp_loops_relevancy_rsc_dat),
      .tile_size_in_rsc_dat(O_tiling_unit_L1_run_cmp_tile_size_in_rsc_dat),
      .tile_size_out_rsc_z(O_tiling_unit_L1_run_cmp_tile_size_out_rsc_z),
      .instr_bound_rsc_z(O_tiling_unit_L1_run_cmp_instr_bound_rsc_z),
      .instr_tile_rsc_z(O_tiling_unit_L1_run_cmp_instr_tile_rsc_z),
      .ccs_ccore_start_rsc_dat(O_tiling_unit_L1_run_cmp_ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(clk),
      .ccs_ccore_srst(rst),
      .ccs_ccore_en(O_tiling_unit_L1_run_cmp_ccs_ccore_en)
    );
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run
      config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3_run_inst
      (
      .clk(clk),
      .rst(rst),
      .layer_instruction_in_rsc_dat(layer_instruction_in_rsc_dat),
      .layer_instruction_in_rsc_vld(layer_instruction_in_rsc_vld),
      .layer_instruction_in_rsc_rdy(layer_instruction_in_rsc_rdy),
      .O_instr_L1_out_rsc_dat(O_instr_L1_out_rsc_dat),
      .O_instr_L1_out_rsc_vld(O_instr_L1_out_rsc_vld),
      .O_instr_L1_out_rsc_rdy(O_instr_L1_out_rsc_rdy),
      .O_instr_L2_out_rsc_dat(O_instr_L2_out_rsc_dat),
      .O_instr_L2_out_rsc_vld(O_instr_L2_out_rsc_vld),
      .O_instr_L2_out_rsc_rdy(O_instr_L2_out_rsc_rdy),
      .O_instr_L3_out_rsc_dat(O_instr_L3_out_rsc_dat),
      .O_instr_L3_out_rsc_vld(O_instr_L3_out_rsc_vld),
      .O_instr_L3_out_rsc_rdy(O_instr_L3_out_rsc_rdy),
      .I_instr_L1_out_rsc_dat(I_instr_L1_out_rsc_dat),
      .I_instr_L1_out_rsc_vld(I_instr_L1_out_rsc_vld),
      .I_instr_L1_out_rsc_rdy(I_instr_L1_out_rsc_rdy),
      .I_instr_L2_out_rsc_dat(I_instr_L2_out_rsc_dat),
      .I_instr_L2_out_rsc_vld(I_instr_L2_out_rsc_vld),
      .I_instr_L2_out_rsc_rdy(I_instr_L2_out_rsc_rdy),
      .I_instr_L3_out_rsc_dat(I_instr_L3_out_rsc_dat),
      .I_instr_L3_out_rsc_vld(I_instr_L3_out_rsc_vld),
      .I_instr_L3_out_rsc_rdy(I_instr_L3_out_rsc_rdy),
      .W_instr_L1_out_rsc_dat(W_instr_L1_out_rsc_dat),
      .W_instr_L1_out_rsc_vld(W_instr_L1_out_rsc_vld),
      .W_instr_L1_out_rsc_rdy(W_instr_L1_out_rsc_rdy),
      .W_instr_L2_out_rsc_dat(W_instr_L2_out_rsc_dat),
      .W_instr_L2_out_rsc_vld(W_instr_L2_out_rsc_vld),
      .W_instr_L2_out_rsc_rdy(W_instr_L2_out_rsc_rdy),
      .W_instr_L3_out_rsc_dat(W_instr_L3_out_rsc_dat),
      .W_instr_L3_out_rsc_vld(W_instr_L3_out_rsc_vld),
      .W_instr_L3_out_rsc_rdy(W_instr_L3_out_rsc_rdy),
      .W_tiling_unit_L3_run_cmp_loops_bound_rsc_dat(W_tiling_unit_L3_run_cmp_loops_bound_rsc_dat),
      .W_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat(W_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat),
      .W_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat(W_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat),
      .W_tiling_unit_L3_run_cmp_instr_bound_rsc_z(W_tiling_unit_L3_run_cmp_instr_bound_rsc_z),
      .W_tiling_unit_L3_run_cmp_instr_tile_rsc_z(W_tiling_unit_L3_run_cmp_instr_tile_rsc_z),
      .W_tiling_unit_L3_run_cmp_ccs_ccore_start_rsc_dat(W_tiling_unit_L3_run_cmp_ccs_ccore_start_rsc_dat),
      .W_tiling_unit_L3_run_cmp_ccs_ccore_en(W_tiling_unit_L3_run_cmp_ccs_ccore_en),
      .ensig_cgo_iro_1(CGHpart_irsig_1),
      .CGHpart_irsig_1(CGHpart_irsig_1),
      .W_tiling_unit_L2_run_cmp_loops_bound_rsc_dat(W_tiling_unit_L2_run_cmp_loops_bound_rsc_dat),
      .W_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat(W_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat),
      .W_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat(W_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat),
      .W_tiling_unit_L2_run_cmp_tile_size_out_rsc_z(W_tiling_unit_L2_run_cmp_tile_size_out_rsc_z),
      .W_tiling_unit_L2_run_cmp_instr_bound_rsc_z(W_tiling_unit_L2_run_cmp_instr_bound_rsc_z),
      .W_tiling_unit_L2_run_cmp_instr_tile_rsc_z(W_tiling_unit_L2_run_cmp_instr_tile_rsc_z),
      .W_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat(W_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat),
      .W_tiling_unit_L2_run_cmp_ccs_ccore_en(W_tiling_unit_L2_run_cmp_ccs_ccore_en),
      .O_tiling_unit_L3_run_cmp_loops_bound_rsc_dat(O_tiling_unit_L3_run_cmp_loops_bound_rsc_dat),
      .O_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat(O_tiling_unit_L3_run_cmp_loops_relevancy_rsc_dat),
      .O_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat(O_tiling_unit_L3_run_cmp_tile_size_in_rsc_dat),
      .O_tiling_unit_L3_run_cmp_instr_bound_rsc_z(O_tiling_unit_L3_run_cmp_instr_bound_rsc_z),
      .O_tiling_unit_L3_run_cmp_instr_tile_rsc_z(O_tiling_unit_L3_run_cmp_instr_tile_rsc_z),
      .O_tiling_unit_L3_run_cmp_ccs_ccore_en(O_tiling_unit_L3_run_cmp_ccs_ccore_en),
      .O_tiling_unit_L2_run_cmp_loops_bound_rsc_dat(O_tiling_unit_L2_run_cmp_loops_bound_rsc_dat),
      .O_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat(O_tiling_unit_L2_run_cmp_loops_relevancy_rsc_dat),
      .O_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat(O_tiling_unit_L2_run_cmp_tile_size_in_rsc_dat),
      .O_tiling_unit_L2_run_cmp_tile_size_out_rsc_z(O_tiling_unit_L2_run_cmp_tile_size_out_rsc_z),
      .O_tiling_unit_L2_run_cmp_instr_bound_rsc_z(O_tiling_unit_L2_run_cmp_instr_bound_rsc_z),
      .O_tiling_unit_L2_run_cmp_instr_tile_rsc_z(O_tiling_unit_L2_run_cmp_instr_tile_rsc_z),
      .O_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat(O_tiling_unit_L2_run_cmp_ccs_ccore_start_rsc_dat),
      .O_tiling_unit_L2_run_cmp_ccs_ccore_en(O_tiling_unit_L2_run_cmp_ccs_ccore_en),
      .O_tiling_unit_L1_run_cmp_loops_bound_rsc_dat(O_tiling_unit_L1_run_cmp_loops_bound_rsc_dat),
      .O_tiling_unit_L1_run_cmp_loops_relevancy_rsc_dat(O_tiling_unit_L1_run_cmp_loops_relevancy_rsc_dat),
      .O_tiling_unit_L1_run_cmp_tile_size_in_rsc_dat(O_tiling_unit_L1_run_cmp_tile_size_in_rsc_dat),
      .O_tiling_unit_L1_run_cmp_tile_size_out_rsc_z(O_tiling_unit_L1_run_cmp_tile_size_out_rsc_z),
      .O_tiling_unit_L1_run_cmp_instr_bound_rsc_z(O_tiling_unit_L1_run_cmp_instr_bound_rsc_z),
      .O_tiling_unit_L1_run_cmp_instr_tile_rsc_z(O_tiling_unit_L1_run_cmp_instr_tile_rsc_z),
      .O_tiling_unit_L1_run_cmp_ccs_ccore_start_rsc_dat(O_tiling_unit_L1_run_cmp_ccs_ccore_start_rsc_dat),
      .O_tiling_unit_L1_run_cmp_ccs_ccore_en(O_tiling_unit_L1_run_cmp_ccs_ccore_en)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1
// ------------------------------------------------------------------


module rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1
    (
  clk, rst, O_wr_data_rsc_dat, O_wr_data_rsc_vld, O_wr_data_rsc_rdy, O_rd_data_rsc_dat,
      O_rd_data_rsc_vld, O_rd_data_rsc_rdy, I_wr_data_rsc_dat, I_wr_data_rsc_vld,
      I_wr_data_rsc_rdy, W_wr_data_rsc_dat, W_wr_data_rsc_vld, W_wr_data_rsc_rdy,
      wr_data_zero_guard_rsc_dat, wr_data_zero_guard_rsc_vld, wr_data_zero_guard_rsc_rdy,
      O_instr_in_rsc_dat, O_instr_in_rsc_vld, O_instr_in_rsc_rdy, I_instr_in_rsc_dat,
      I_instr_in_rsc_vld, I_instr_in_rsc_rdy, W_instr_in_rsc_dat, W_instr_in_rsc_vld,
      W_instr_in_rsc_rdy
);
  input clk;
  input rst;
  input [15:0] O_wr_data_rsc_dat;
  input O_wr_data_rsc_vld;
  output O_wr_data_rsc_rdy;
  output [15:0] O_rd_data_rsc_dat;
  output O_rd_data_rsc_vld;
  input O_rd_data_rsc_rdy;
  input [15:0] I_wr_data_rsc_dat;
  input I_wr_data_rsc_vld;
  output I_wr_data_rsc_rdy;
  input [15:0] W_wr_data_rsc_dat;
  input W_wr_data_rsc_vld;
  output W_wr_data_rsc_rdy;
  input wr_data_zero_guard_rsc_dat;
  input wr_data_zero_guard_rsc_vld;
  output wr_data_zero_guard_rsc_rdy;
  input [49:0] O_instr_in_rsc_dat;
  input O_instr_in_rsc_vld;
  output O_instr_in_rsc_rdy;
  input [49:0] I_instr_in_rsc_dat;
  input I_instr_in_rsc_vld;
  output I_instr_in_rsc_rdy;
  input [49:0] W_instr_in_rsc_dat;
  input W_instr_in_rsc_vld;
  output W_instr_in_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run
      rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1_run_inst
      (
      .clk(clk),
      .rst(rst),
      .O_wr_data_rsc_dat(O_wr_data_rsc_dat),
      .O_wr_data_rsc_vld(O_wr_data_rsc_vld),
      .O_wr_data_rsc_rdy(O_wr_data_rsc_rdy),
      .O_rd_data_rsc_dat(O_rd_data_rsc_dat),
      .O_rd_data_rsc_vld(O_rd_data_rsc_vld),
      .O_rd_data_rsc_rdy(O_rd_data_rsc_rdy),
      .I_wr_data_rsc_dat(I_wr_data_rsc_dat),
      .I_wr_data_rsc_vld(I_wr_data_rsc_vld),
      .I_wr_data_rsc_rdy(I_wr_data_rsc_rdy),
      .W_wr_data_rsc_dat(W_wr_data_rsc_dat),
      .W_wr_data_rsc_vld(W_wr_data_rsc_vld),
      .W_wr_data_rsc_rdy(W_wr_data_rsc_rdy),
      .wr_data_zero_guard_rsc_dat(wr_data_zero_guard_rsc_dat),
      .wr_data_zero_guard_rsc_vld(wr_data_zero_guard_rsc_vld),
      .wr_data_zero_guard_rsc_rdy(wr_data_zero_guard_rsc_rdy),
      .O_instr_in_rsc_dat(O_instr_in_rsc_dat),
      .O_instr_in_rsc_vld(O_instr_in_rsc_vld),
      .O_instr_in_rsc_rdy(O_instr_in_rsc_rdy),
      .I_instr_in_rsc_dat(I_instr_in_rsc_dat),
      .I_instr_in_rsc_vld(I_instr_in_rsc_vld),
      .I_instr_in_rsc_rdy(I_instr_in_rsc_rdy),
      .W_instr_in_rsc_dat(W_instr_in_rsc_dat),
      .W_instr_in_rsc_vld(W_instr_in_rsc_vld),
      .W_instr_in_rsc_rdy(W_instr_in_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_partial_000001
// ------------------------------------------------------------------


module top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_partial_000001
    (
  clk, rst, O_data_in_rsc_dat_data, O_data_in_rsc_vld, O_data_in_rsc_rdy, O_data_out_rsc_dat_data,
      O_data_out_rsc_vld, O_data_out_rsc_rdy, I_data_in_rsc_dat_data, I_data_in_rsc_vld,
      I_data_in_rsc_rdy, W_data_in_rsc_dat_data, W_data_in_rsc_vld, W_data_in_rsc_rdy,
      zero_guard_in_rsc_dat, zero_guard_in_rsc_vld, zero_guard_in_rsc_rdy, layer_instruction_in_rsc_dat_relevancy,
      layer_instruction_in_rsc_dat_bound, layer_instruction_in_rsc_dat_relevancy_1,
      layer_instruction_in_rsc_dat_bound_1, layer_instruction_in_rsc_dat_relevancy_2,
      layer_instruction_in_rsc_dat_bound_2, layer_instruction_in_rsc_dat_relevancy_3,
      layer_instruction_in_rsc_dat_bound_3, layer_instruction_in_rsc_dat_relevancy_4,
      layer_instruction_in_rsc_dat_bound_4, layer_instruction_in_rsc_dat_relevancy_5,
      layer_instruction_in_rsc_dat_bound_5, layer_instruction_in_rsc_dat_relevancy_6,
      layer_instruction_in_rsc_dat_bound_6, layer_instruction_in_rsc_dat_relevancy_7,
      layer_instruction_in_rsc_dat_bound_7, layer_instruction_in_rsc_dat_relevancy_8,
      layer_instruction_in_rsc_dat_bound_8, layer_instruction_in_rsc_vld, layer_instruction_in_rsc_rdy
);
  input clk;
  input rst;
  input [15:0] O_data_in_rsc_dat_data;
  input O_data_in_rsc_vld;
  output O_data_in_rsc_rdy;
  output [15:0] O_data_out_rsc_dat_data;
  output O_data_out_rsc_vld;
  input O_data_out_rsc_rdy;
  input [15:0] I_data_in_rsc_dat_data;
  input I_data_in_rsc_vld;
  output I_data_in_rsc_rdy;
  input [15:0] W_data_in_rsc_dat_data;
  input W_data_in_rsc_vld;
  output W_data_in_rsc_rdy;
  input zero_guard_in_rsc_dat;
  input zero_guard_in_rsc_vld;
  output zero_guard_in_rsc_rdy;
  input [4:0] layer_instruction_in_rsc_dat_relevancy;
  input [24:0] layer_instruction_in_rsc_dat_bound;
  input [4:0] layer_instruction_in_rsc_dat_relevancy_1;
  input [54:0] layer_instruction_in_rsc_dat_bound_1;
  input [4:0] layer_instruction_in_rsc_dat_relevancy_2;
  input [79:0] layer_instruction_in_rsc_dat_bound_2;
  input [4:0] layer_instruction_in_rsc_dat_relevancy_3;
  input [24:0] layer_instruction_in_rsc_dat_bound_3;
  input [4:0] layer_instruction_in_rsc_dat_relevancy_4;
  input [44:0] layer_instruction_in_rsc_dat_bound_4;
  input [4:0] layer_instruction_in_rsc_dat_relevancy_5;
  input [69:0] layer_instruction_in_rsc_dat_bound_5;
  input [4:0] layer_instruction_in_rsc_dat_relevancy_6;
  input [24:0] layer_instruction_in_rsc_dat_bound_6;
  input [4:0] layer_instruction_in_rsc_dat_relevancy_7;
  input [44:0] layer_instruction_in_rsc_dat_bound_7;
  input [4:0] layer_instruction_in_rsc_dat_relevancy_8;
  input [69:0] layer_instruction_in_rsc_dat_bound_8;
  input layer_instruction_in_rsc_vld;
  output layer_instruction_in_rsc_rdy;


  // Interconnect Declarations
  wire [49:0] O_instr_L1_out_rsc_dat_nCCInst;
  wire [89:0] O_instr_L2_out_rsc_dat_nCCInst;
  wire [139:0] O_instr_L3_out_rsc_dat_nCCInst;
  wire [49:0] I_instr_L1_out_rsc_dat_nCCInst;
  wire [89:0] I_instr_L2_out_rsc_dat_nCCInst;
  wire [139:0] I_instr_L3_out_rsc_dat_nCCInst;
  wire [49:0] W_instr_L1_out_rsc_dat_nCCInst;
  wire [109:0] W_instr_L2_out_rsc_dat_nCCInst;
  wire [159:0] W_instr_L3_out_rsc_dat_nCCInst;
  wire [15:0] O_rd_data_rsc_dat_nPE;
  wire layer_instruction_in_rsc_rdy_nCCInst_bud;
  wire O_instr_L1_out_rsc_vld_nCCInst_bud;
  wire O_instr_in_rsc_rdy_nPE_bud;
  wire O_instr_L2_out_rsc_vld_nCCInst_bud;
  wire O_instr_L3_out_rsc_vld_nCCInst_bud;
  wire I_instr_L1_out_rsc_vld_nCCInst_bud;
  wire I_instr_in_rsc_rdy_nPE_bud;
  wire I_instr_L2_out_rsc_vld_nCCInst_bud;
  wire I_instr_L3_out_rsc_vld_nCCInst_bud;
  wire W_instr_L1_out_rsc_vld_nCCInst_bud;
  wire W_instr_in_rsc_rdy_nPE_bud;
  wire W_instr_L2_out_rsc_vld_nCCInst_bud;
  wire W_instr_L3_out_rsc_vld_nCCInst_bud;
  wire O_wr_data_rsc_rdy_nPE_bud;
  wire O_rd_data_rsc_vld_nPE_bud;
  wire I_wr_data_rsc_rdy_nPE_bud;
  wire W_wr_data_rsc_rdy_nPE_bud;
  wire wr_data_zero_guard_rsc_rdy_nPE_bud;


  // Interconnect Declarations for Component Instantiations 
  wire [484:0] nl_CCInst_layer_instruction_in_rsc_dat;
  assign nl_CCInst_layer_instruction_in_rsc_dat = {layer_instruction_in_rsc_dat_relevancy
      , layer_instruction_in_rsc_dat_bound , layer_instruction_in_rsc_dat_relevancy_1
      , layer_instruction_in_rsc_dat_bound_1 , layer_instruction_in_rsc_dat_relevancy_2
      , layer_instruction_in_rsc_dat_bound_2 , layer_instruction_in_rsc_dat_relevancy_3
      , layer_instruction_in_rsc_dat_bound_3 , layer_instruction_in_rsc_dat_relevancy_4
      , layer_instruction_in_rsc_dat_bound_4 , layer_instruction_in_rsc_dat_relevancy_5
      , layer_instruction_in_rsc_dat_bound_5 , layer_instruction_in_rsc_dat_relevancy_6
      , layer_instruction_in_rsc_dat_bound_6 , layer_instruction_in_rsc_dat_relevancy_7
      , layer_instruction_in_rsc_dat_bound_7 , layer_instruction_in_rsc_dat_relevancy_8
      , layer_instruction_in_rsc_dat_bound_8};
  config_control_unit_5_O_addr_type_L1_O_addr_type_L2_O_addr_type_L3_I_addr_type_L1_I_addr_type_L2_I_addr_type_L3_W_addr_type_L1_W_addr_type_L2_W_addr_type_L3
      CCInst (
      .clk(clk),
      .rst(rst),
      .layer_instruction_in_rsc_dat(nl_CCInst_layer_instruction_in_rsc_dat[484:0]),
      .layer_instruction_in_rsc_vld(layer_instruction_in_rsc_vld),
      .layer_instruction_in_rsc_rdy(layer_instruction_in_rsc_rdy_nCCInst_bud),
      .O_instr_L1_out_rsc_dat(O_instr_L1_out_rsc_dat_nCCInst),
      .O_instr_L1_out_rsc_vld(O_instr_L1_out_rsc_vld_nCCInst_bud),
      .O_instr_L1_out_rsc_rdy(O_instr_in_rsc_rdy_nPE_bud),
      .O_instr_L2_out_rsc_dat(O_instr_L2_out_rsc_dat_nCCInst),
      .O_instr_L2_out_rsc_vld(O_instr_L2_out_rsc_vld_nCCInst_bud),
      .O_instr_L2_out_rsc_rdy(1'b1),
      .O_instr_L3_out_rsc_dat(O_instr_L3_out_rsc_dat_nCCInst),
      .O_instr_L3_out_rsc_vld(O_instr_L3_out_rsc_vld_nCCInst_bud),
      .O_instr_L3_out_rsc_rdy(1'b1),
      .I_instr_L1_out_rsc_dat(I_instr_L1_out_rsc_dat_nCCInst),
      .I_instr_L1_out_rsc_vld(I_instr_L1_out_rsc_vld_nCCInst_bud),
      .I_instr_L1_out_rsc_rdy(I_instr_in_rsc_rdy_nPE_bud),
      .I_instr_L2_out_rsc_dat(I_instr_L2_out_rsc_dat_nCCInst),
      .I_instr_L2_out_rsc_vld(I_instr_L2_out_rsc_vld_nCCInst_bud),
      .I_instr_L2_out_rsc_rdy(1'b1),
      .I_instr_L3_out_rsc_dat(I_instr_L3_out_rsc_dat_nCCInst),
      .I_instr_L3_out_rsc_vld(I_instr_L3_out_rsc_vld_nCCInst_bud),
      .I_instr_L3_out_rsc_rdy(1'b1),
      .W_instr_L1_out_rsc_dat(W_instr_L1_out_rsc_dat_nCCInst),
      .W_instr_L1_out_rsc_vld(W_instr_L1_out_rsc_vld_nCCInst_bud),
      .W_instr_L1_out_rsc_rdy(W_instr_in_rsc_rdy_nPE_bud),
      .W_instr_L2_out_rsc_dat(W_instr_L2_out_rsc_dat_nCCInst),
      .W_instr_L2_out_rsc_vld(W_instr_L2_out_rsc_vld_nCCInst_bud),
      .W_instr_L2_out_rsc_rdy(1'b1),
      .W_instr_L3_out_rsc_dat(W_instr_L3_out_rsc_dat_nCCInst),
      .W_instr_L3_out_rsc_vld(W_instr_L3_out_rsc_vld_nCCInst_bud),
      .W_instr_L3_out_rsc_rdy(1'b1)
    );
  rf_5_32_32_32_1_1_1_1_1_1_O_partial_type_O_addr_type_L1_I_type_I_addr_type_L1_W_type_W_addr_type_L1
      PE (
      .clk(clk),
      .rst(rst),
      .O_wr_data_rsc_dat(O_data_in_rsc_dat_data),
      .O_wr_data_rsc_vld(O_data_in_rsc_vld),
      .O_wr_data_rsc_rdy(O_wr_data_rsc_rdy_nPE_bud),
      .O_rd_data_rsc_dat(O_rd_data_rsc_dat_nPE),
      .O_rd_data_rsc_vld(O_rd_data_rsc_vld_nPE_bud),
      .O_rd_data_rsc_rdy(O_data_out_rsc_rdy),
      .I_wr_data_rsc_dat(I_data_in_rsc_dat_data),
      .I_wr_data_rsc_vld(I_data_in_rsc_vld),
      .I_wr_data_rsc_rdy(I_wr_data_rsc_rdy_nPE_bud),
      .W_wr_data_rsc_dat(W_data_in_rsc_dat_data),
      .W_wr_data_rsc_vld(W_data_in_rsc_vld),
      .W_wr_data_rsc_rdy(W_wr_data_rsc_rdy_nPE_bud),
      .wr_data_zero_guard_rsc_dat(zero_guard_in_rsc_dat),
      .wr_data_zero_guard_rsc_vld(zero_guard_in_rsc_vld),
      .wr_data_zero_guard_rsc_rdy(wr_data_zero_guard_rsc_rdy_nPE_bud),
      .O_instr_in_rsc_dat(O_instr_L1_out_rsc_dat_nCCInst),
      .O_instr_in_rsc_vld(O_instr_L1_out_rsc_vld_nCCInst_bud),
      .O_instr_in_rsc_rdy(O_instr_in_rsc_rdy_nPE_bud),
      .I_instr_in_rsc_dat(I_instr_L1_out_rsc_dat_nCCInst),
      .I_instr_in_rsc_vld(I_instr_L1_out_rsc_vld_nCCInst_bud),
      .I_instr_in_rsc_rdy(I_instr_in_rsc_rdy_nPE_bud),
      .W_instr_in_rsc_dat(W_instr_L1_out_rsc_dat_nCCInst),
      .W_instr_in_rsc_vld(W_instr_L1_out_rsc_vld_nCCInst_bud),
      .W_instr_in_rsc_rdy(W_instr_in_rsc_rdy_nPE_bud)
    );
  assign O_data_out_rsc_dat_data = O_rd_data_rsc_dat_nPE;
  assign layer_instruction_in_rsc_rdy = layer_instruction_in_rsc_rdy_nCCInst_bud;
  assign O_data_in_rsc_rdy = O_wr_data_rsc_rdy_nPE_bud;
  assign O_data_out_rsc_vld = O_rd_data_rsc_vld_nPE_bud;
  assign I_data_in_rsc_rdy = I_wr_data_rsc_rdy_nPE_bud;
  assign W_data_in_rsc_rdy = W_wr_data_rsc_rdy_nPE_bud;
  assign zero_guard_in_rsc_rdy = wr_data_zero_guard_rsc_rdy_nPE_bud;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_partial_000000
// ------------------------------------------------------------------


module top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_partial_000000
    (
  clk, rst, O_data_in_rsc_dat, O_data_in_rsc_vld, O_data_in_rsc_rdy, O_data_out_rsc_dat,
      O_data_out_rsc_vld, O_data_out_rsc_rdy, I_data_in_rsc_dat, I_data_in_rsc_vld,
      I_data_in_rsc_rdy, W_data_in_rsc_dat, W_data_in_rsc_vld, W_data_in_rsc_rdy,
      zero_guard_in_rsc_dat, zero_guard_in_rsc_vld, zero_guard_in_rsc_rdy, layer_instruction_in_rsc_dat,
      layer_instruction_in_rsc_vld, layer_instruction_in_rsc_rdy
);
  input clk;
  input rst;
  input [15:0] O_data_in_rsc_dat;
  input O_data_in_rsc_vld;
  output O_data_in_rsc_rdy;
  output [15:0] O_data_out_rsc_dat;
  output O_data_out_rsc_vld;
  input O_data_out_rsc_rdy;
  input [15:0] I_data_in_rsc_dat;
  input I_data_in_rsc_vld;
  output I_data_in_rsc_rdy;
  input [15:0] W_data_in_rsc_dat;
  input W_data_in_rsc_vld;
  output W_data_in_rsc_rdy;
  input zero_guard_in_rsc_dat;
  input zero_guard_in_rsc_vld;
  output zero_guard_in_rsc_rdy;
  input [484:0] layer_instruction_in_rsc_dat;
  input layer_instruction_in_rsc_vld;
  output layer_instruction_in_rsc_rdy;


  // Interconnect Declarations
  wire [15:0] O_data_out_rsc_dat_data;


  // Interconnect Declarations for Component Instantiations 
  wire [4:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000000;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000000
      = layer_instruction_in_rsc_dat[484:480];
  wire [24:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000001;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000001
      = layer_instruction_in_rsc_dat[479:455];
  wire [4:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000002;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000002
      = layer_instruction_in_rsc_dat[454:450];
  wire [54:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000003;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000003
      = layer_instruction_in_rsc_dat[449:395];
  wire [4:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000004;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000004
      = layer_instruction_in_rsc_dat[394:390];
  wire [79:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000005;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000005
      = layer_instruction_in_rsc_dat[389:310];
  wire [4:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000006;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000006
      = layer_instruction_in_rsc_dat[309:305];
  wire [24:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000007;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000007
      = layer_instruction_in_rsc_dat[304:280];
  wire [4:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000008;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000008
      = layer_instruction_in_rsc_dat[279:275];
  wire [44:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000009;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000009
      = layer_instruction_in_rsc_dat[274:230];
  wire [4:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000010;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000010
      = layer_instruction_in_rsc_dat[229:225];
  wire [69:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000011;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000011
      = layer_instruction_in_rsc_dat[224:155];
  wire [4:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000012;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000012
      = layer_instruction_in_rsc_dat[154:150];
  wire [24:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000013;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000013
      = layer_instruction_in_rsc_dat[149:125];
  wire [4:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000014;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000014
      = layer_instruction_in_rsc_dat[124:120];
  wire [44:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000015;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000015
      = layer_instruction_in_rsc_dat[119:75];
  wire [4:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000016;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000016
      = layer_instruction_in_rsc_dat[74:70];
  wire [69:0] nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000017;
  assign nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000017
      = layer_instruction_in_rsc_dat[69:0];
  top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_partial_000001
      top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_partial_000002
      (
      .clk(clk),
      .rst(rst),
      .O_data_in_rsc_dat_data(O_data_in_rsc_dat),
      .O_data_in_rsc_vld(O_data_in_rsc_vld),
      .O_data_in_rsc_rdy(O_data_in_rsc_rdy),
      .O_data_out_rsc_dat_data(O_data_out_rsc_dat_data),
      .O_data_out_rsc_vld(O_data_out_rsc_vld),
      .O_data_out_rsc_rdy(O_data_out_rsc_rdy),
      .I_data_in_rsc_dat_data(I_data_in_rsc_dat),
      .I_data_in_rsc_vld(I_data_in_rsc_vld),
      .I_data_in_rsc_rdy(I_data_in_rsc_rdy),
      .W_data_in_rsc_dat_data(W_data_in_rsc_dat),
      .W_data_in_rsc_vld(W_data_in_rsc_vld),
      .W_data_in_rsc_rdy(W_data_in_rsc_rdy),
      .zero_guard_in_rsc_dat(zero_guard_in_rsc_dat),
      .zero_guard_in_rsc_vld(zero_guard_in_rsc_vld),
      .zero_guard_in_rsc_rdy(zero_guard_in_rsc_rdy),
      .layer_instruction_in_rsc_dat_relevancy(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000000[4:0]),
      .layer_instruction_in_rsc_dat_bound(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000001[24:0]),
      .layer_instruction_in_rsc_dat_relevancy_1(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000002[4:0]),
      .layer_instruction_in_rsc_dat_bound_1(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000003[54:0]),
      .layer_instruction_in_rsc_dat_relevancy_2(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000004[4:0]),
      .layer_instruction_in_rsc_dat_bound_2(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000005[79:0]),
      .layer_instruction_in_rsc_dat_relevancy_3(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000006[4:0]),
      .layer_instruction_in_rsc_dat_bound_3(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000007[24:0]),
      .layer_instruction_in_rsc_dat_relevancy_4(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000008[4:0]),
      .layer_instruction_in_rsc_dat_bound_4(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000009[44:0]),
      .layer_instruction_in_rsc_dat_relevancy_5(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000010[4:0]),
      .layer_instruction_in_rsc_dat_bound_5(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000011[69:0]),
      .layer_instruction_in_rsc_dat_relevancy_6(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000012[4:0]),
      .layer_instruction_in_rsc_dat_bound_6(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000013[24:0]),
      .layer_instruction_in_rsc_dat_relevancy_7(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000014[4:0]),
      .layer_instruction_in_rsc_dat_bound_7(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000015[44:0]),
      .layer_instruction_in_rsc_dat_relevancy_8(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000016[4:0]),
      .layer_instruction_in_rsc_dat_bound_8(nl_top_5_32_1_1_O_addr_type_L1_32_1_1_I_addr_type_L1_32_1_1_W_addr_type_L1_5_288_8_8_O_addr_type_L2_312_8_8_I_addr_type_L2_1728_8_8_W_addr_type_L2_5_8640_8_8_O_addr_type_L3_8640_8_8_I_addr_type_L3_55296_8_8_W_addr_type_L3_O_parti000017[69:0]),
      .layer_instruction_in_rsc_vld(layer_instruction_in_rsc_vld),
      .layer_instruction_in_rsc_rdy(layer_instruction_in_rsc_rdy)
    );
  assign O_data_out_rsc_dat = O_data_out_rsc_dat_data;
endmodule



